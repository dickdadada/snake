module rom_snakeg (clock, address, q);
input clock;
output [7:0] q;
input [11:0] address;
reg [7:0] dout;
reg [7:0] ram [4095:0];
assign q = dout;

initial begin
  ram[0]  = 128;
  ram[1]  = 133;
  ram[2]  = 130;
  ram[3]  = 130;
  ram[4]  = 129;
  ram[5]  = 127;
  ram[6]  = 129;
  ram[7]  = 129;
  ram[8]  = 128;
  ram[9]  = 128;
  ram[10]  = 128;
  ram[11]  = 128;
  ram[12]  = 129;
  ram[13]  = 129;
  ram[14]  = 129;
  ram[15]  = 129;
  ram[16]  = 130;
  ram[17]  = 130;
  ram[18]  = 130;
  ram[19]  = 130;
  ram[20]  = 130;
  ram[21]  = 130;
  ram[22]  = 130;
  ram[23]  = 130;
  ram[24]  = 130;
  ram[25]  = 130;
  ram[26]  = 130;
  ram[27]  = 130;
  ram[28]  = 130;
  ram[29]  = 130;
  ram[30]  = 130;
  ram[31]  = 130;
  ram[32]  = 130;
  ram[33]  = 130;
  ram[34]  = 130;
  ram[35]  = 130;
  ram[36]  = 130;
  ram[37]  = 130;
  ram[38]  = 130;
  ram[39]  = 130;
  ram[40]  = 130;
  ram[41]  = 130;
  ram[42]  = 130;
  ram[43]  = 130;
  ram[44]  = 130;
  ram[45]  = 130;
  ram[46]  = 130;
  ram[47]  = 130;
  ram[48]  = 130;
  ram[49]  = 130;
  ram[50]  = 129;
  ram[51]  = 129;
  ram[52]  = 129;
  ram[53]  = 129;
  ram[54]  = 129;
  ram[55]  = 129;
  ram[56]  = 128;
  ram[57]  = 129;
  ram[58]  = 129;
  ram[59]  = 129;
  ram[60]  = 129;
  ram[61]  = 129;
  ram[62]  = 129;
  ram[63]  = 127;
  ram[64]  = 131;
  ram[65]  = 135;
  ram[66]  = 132;
  ram[67]  = 132;
  ram[68]  = 132;
  ram[69]  = 130;
  ram[70]  = 132;
  ram[71]  = 131;
  ram[72]  = 131;
  ram[73]  = 131;
  ram[74]  = 131;
  ram[75]  = 131;
  ram[76]  = 132;
  ram[77]  = 132;
  ram[78]  = 132;
  ram[79]  = 132;
  ram[80]  = 132;
  ram[81]  = 132;
  ram[82]  = 132;
  ram[83]  = 132;
  ram[84]  = 132;
  ram[85]  = 132;
  ram[86]  = 132;
  ram[87]  = 132;
  ram[88]  = 132;
  ram[89]  = 132;
  ram[90]  = 132;
  ram[91]  = 132;
  ram[92]  = 132;
  ram[93]  = 132;
  ram[94]  = 132;
  ram[95]  = 132;
  ram[96]  = 132;
  ram[97]  = 132;
  ram[98]  = 132;
  ram[99]  = 132;
  ram[100]  = 132;
  ram[101]  = 132;
  ram[102]  = 132;
  ram[103]  = 132;
  ram[104]  = 132;
  ram[105]  = 132;
  ram[106]  = 132;
  ram[107]  = 132;
  ram[108]  = 132;
  ram[109]  = 132;
  ram[110]  = 132;
  ram[111]  = 132;
  ram[112]  = 132;
  ram[113]  = 132;
  ram[114]  = 131;
  ram[115]  = 131;
  ram[116]  = 131;
  ram[117]  = 131;
  ram[118]  = 131;
  ram[119]  = 131;
  ram[120]  = 131;
  ram[121]  = 131;
  ram[122]  = 131;
  ram[123]  = 131;
  ram[124]  = 132;
  ram[125]  = 132;
  ram[126]  = 132;
  ram[127]  = 129;
  ram[128]  = 132;
  ram[129]  = 136;
  ram[130]  = 131;
  ram[131]  = 132;
  ram[132]  = 133;
  ram[133]  = 132;
  ram[134]  = 132;
  ram[135]  = 132;
  ram[136]  = 133;
  ram[137]  = 133;
  ram[138]  = 132;
  ram[139]  = 132;
  ram[140]  = 132;
  ram[141]  = 132;
  ram[142]  = 133;
  ram[143]  = 133;
  ram[144]  = 132;
  ram[145]  = 132;
  ram[146]  = 132;
  ram[147]  = 132;
  ram[148]  = 132;
  ram[149]  = 132;
  ram[150]  = 132;
  ram[151]  = 132;
  ram[152]  = 132;
  ram[153]  = 132;
  ram[154]  = 132;
  ram[155]  = 132;
  ram[156]  = 132;
  ram[157]  = 132;
  ram[158]  = 132;
  ram[159]  = 132;
  ram[160]  = 132;
  ram[161]  = 132;
  ram[162]  = 132;
  ram[163]  = 132;
  ram[164]  = 132;
  ram[165]  = 132;
  ram[166]  = 132;
  ram[167]  = 132;
  ram[168]  = 132;
  ram[169]  = 132;
  ram[170]  = 132;
  ram[171]  = 132;
  ram[172]  = 132;
  ram[173]  = 132;
  ram[174]  = 132;
  ram[175]  = 132;
  ram[176]  = 133;
  ram[177]  = 133;
  ram[178]  = 132;
  ram[179]  = 132;
  ram[180]  = 132;
  ram[181]  = 132;
  ram[182]  = 132;
  ram[183]  = 132;
  ram[184]  = 132;
  ram[185]  = 132;
  ram[186]  = 132;
  ram[187]  = 132;
  ram[188]  = 132;
  ram[189]  = 133;
  ram[190]  = 132;
  ram[191]  = 130;
  ram[192]  = 132;
  ram[193]  = 135;
  ram[194]  = 130;
  ram[195]  = 131;
  ram[196]  = 133;
  ram[197]  = 132;
  ram[198]  = 132;
  ram[199]  = 131;
  ram[200]  = 133;
  ram[201]  = 133;
  ram[202]  = 133;
  ram[203]  = 133;
  ram[204]  = 133;
  ram[205]  = 133;
  ram[206]  = 134;
  ram[207]  = 134;
  ram[208]  = 132;
  ram[209]  = 132;
  ram[210]  = 132;
  ram[211]  = 132;
  ram[212]  = 132;
  ram[213]  = 132;
  ram[214]  = 132;
  ram[215]  = 132;
  ram[216]  = 132;
  ram[217]  = 132;
  ram[218]  = 132;
  ram[219]  = 132;
  ram[220]  = 132;
  ram[221]  = 132;
  ram[222]  = 132;
  ram[223]  = 132;
  ram[224]  = 132;
  ram[225]  = 132;
  ram[226]  = 132;
  ram[227]  = 132;
  ram[228]  = 132;
  ram[229]  = 132;
  ram[230]  = 132;
  ram[231]  = 132;
  ram[232]  = 132;
  ram[233]  = 132;
  ram[234]  = 132;
  ram[235]  = 132;
  ram[236]  = 132;
  ram[237]  = 132;
  ram[238]  = 132;
  ram[239]  = 132;
  ram[240]  = 133;
  ram[241]  = 133;
  ram[242]  = 132;
  ram[243]  = 132;
  ram[244]  = 132;
  ram[245]  = 132;
  ram[246]  = 132;
  ram[247]  = 132;
  ram[248]  = 131;
  ram[249]  = 132;
  ram[250]  = 132;
  ram[251]  = 131;
  ram[252]  = 132;
  ram[253]  = 132;
  ram[254]  = 132;
  ram[255]  = 130;
  ram[256]  = 132;
  ram[257]  = 136;
  ram[258]  = 131;
  ram[259]  = 131;
  ram[260]  = 133;
  ram[261]  = 132;
  ram[262]  = 131;
  ram[263]  = 130;
  ram[264]  = 133;
  ram[265]  = 133;
  ram[266]  = 133;
  ram[267]  = 133;
  ram[268]  = 133;
  ram[269]  = 133;
  ram[270]  = 133;
  ram[271]  = 133;
  ram[272]  = 133;
  ram[273]  = 133;
  ram[274]  = 133;
  ram[275]  = 133;
  ram[276]  = 132;
  ram[277]  = 132;
  ram[278]  = 132;
  ram[279]  = 132;
  ram[280]  = 132;
  ram[281]  = 132;
  ram[282]  = 132;
  ram[283]  = 132;
  ram[284]  = 133;
  ram[285]  = 133;
  ram[286]  = 133;
  ram[287]  = 133;
  ram[288]  = 133;
  ram[289]  = 133;
  ram[290]  = 133;
  ram[291]  = 133;
  ram[292]  = 133;
  ram[293]  = 133;
  ram[294]  = 133;
  ram[295]  = 133;
  ram[296]  = 133;
  ram[297]  = 133;
  ram[298]  = 133;
  ram[299]  = 133;
  ram[300]  = 133;
  ram[301]  = 133;
  ram[302]  = 133;
  ram[303]  = 133;
  ram[304]  = 133;
  ram[305]  = 133;
  ram[306]  = 133;
  ram[307]  = 133;
  ram[308]  = 133;
  ram[309]  = 133;
  ram[310]  = 133;
  ram[311]  = 133;
  ram[312]  = 132;
  ram[313]  = 132;
  ram[314]  = 132;
  ram[315]  = 132;
  ram[316]  = 132;
  ram[317]  = 133;
  ram[318]  = 131;
  ram[319]  = 129;
  ram[320]  = 132;
  ram[321]  = 136;
  ram[322]  = 131;
  ram[323]  = 131;
  ram[324]  = 133;
  ram[325]  = 131;
  ram[326]  = 131;
  ram[327]  = 130;
  ram[328]  = 132;
  ram[329]  = 132;
  ram[330]  = 132;
  ram[331]  = 132;
  ram[332]  = 131;
  ram[333]  = 132;
  ram[334]  = 132;
  ram[335]  = 132;
  ram[336]  = 132;
  ram[337]  = 132;
  ram[338]  = 132;
  ram[339]  = 132;
  ram[340]  = 131;
  ram[341]  = 131;
  ram[342]  = 131;
  ram[343]  = 131;
  ram[344]  = 131;
  ram[345]  = 131;
  ram[346]  = 131;
  ram[347]  = 131;
  ram[348]  = 132;
  ram[349]  = 132;
  ram[350]  = 132;
  ram[351]  = 132;
  ram[352]  = 132;
  ram[353]  = 132;
  ram[354]  = 132;
  ram[355]  = 132;
  ram[356]  = 132;
  ram[357]  = 132;
  ram[358]  = 132;
  ram[359]  = 132;
  ram[360]  = 132;
  ram[361]  = 132;
  ram[362]  = 132;
  ram[363]  = 132;
  ram[364]  = 132;
  ram[365]  = 132;
  ram[366]  = 132;
  ram[367]  = 132;
  ram[368]  = 132;
  ram[369]  = 132;
  ram[370]  = 132;
  ram[371]  = 132;
  ram[372]  = 132;
  ram[373]  = 132;
  ram[374]  = 132;
  ram[375]  = 132;
  ram[376]  = 132;
  ram[377]  = 132;
  ram[378]  = 132;
  ram[379]  = 132;
  ram[380]  = 132;
  ram[381]  = 132;
  ram[382]  = 131;
  ram[383]  = 129;
  ram[384]  = 130;
  ram[385]  = 134;
  ram[386]  = 131;
  ram[387]  = 131;
  ram[388]  = 131;
  ram[389]  = 130;
  ram[390]  = 131;
  ram[391]  = 130;
  ram[392]  = 131;
  ram[393]  = 131;
  ram[394]  = 131;
  ram[395]  = 131;
  ram[396]  = 130;
  ram[397]  = 130;
  ram[398]  = 130;
  ram[399]  = 130;
  ram[400]  = 131;
  ram[401]  = 131;
  ram[402]  = 131;
  ram[403]  = 131;
  ram[404]  = 130;
  ram[405]  = 130;
  ram[406]  = 130;
  ram[407]  = 130;
  ram[408]  = 130;
  ram[409]  = 130;
  ram[410]  = 130;
  ram[411]  = 130;
  ram[412]  = 130;
  ram[413]  = 130;
  ram[414]  = 130;
  ram[415]  = 130;
  ram[416]  = 130;
  ram[417]  = 130;
  ram[418]  = 130;
  ram[419]  = 130;
  ram[420]  = 130;
  ram[421]  = 130;
  ram[422]  = 130;
  ram[423]  = 130;
  ram[424]  = 130;
  ram[425]  = 130;
  ram[426]  = 130;
  ram[427]  = 130;
  ram[428]  = 131;
  ram[429]  = 131;
  ram[430]  = 131;
  ram[431]  = 131;
  ram[432]  = 131;
  ram[433]  = 131;
  ram[434]  = 131;
  ram[435]  = 131;
  ram[436]  = 130;
  ram[437]  = 130;
  ram[438]  = 130;
  ram[439]  = 130;
  ram[440]  = 131;
  ram[441]  = 131;
  ram[442]  = 131;
  ram[443]  = 130;
  ram[444]  = 132;
  ram[445]  = 132;
  ram[446]  = 130;
  ram[447]  = 128;
  ram[448]  = 130;
  ram[449]  = 135;
  ram[450]  = 132;
  ram[451]  = 132;
  ram[452]  = 132;
  ram[453]  = 130;
  ram[454]  = 131;
  ram[455]  = 132;
  ram[456]  = 132;
  ram[457]  = 133;
  ram[458]  = 132;
  ram[459]  = 132;
  ram[460]  = 131;
  ram[461]  = 131;
  ram[462]  = 131;
  ram[463]  = 131;
  ram[464]  = 131;
  ram[465]  = 132;
  ram[466]  = 132;
  ram[467]  = 132;
  ram[468]  = 131;
  ram[469]  = 131;
  ram[470]  = 131;
  ram[471]  = 131;
  ram[472]  = 131;
  ram[473]  = 131;
  ram[474]  = 131;
  ram[475]  = 131;
  ram[476]  = 131;
  ram[477]  = 131;
  ram[478]  = 131;
  ram[479]  = 131;
  ram[480]  = 131;
  ram[481]  = 131;
  ram[482]  = 131;
  ram[483]  = 131;
  ram[484]  = 131;
  ram[485]  = 131;
  ram[486]  = 131;
  ram[487]  = 131;
  ram[488]  = 131;
  ram[489]  = 131;
  ram[490]  = 131;
  ram[491]  = 131;
  ram[492]  = 132;
  ram[493]  = 132;
  ram[494]  = 132;
  ram[495]  = 132;
  ram[496]  = 132;
  ram[497]  = 132;
  ram[498]  = 132;
  ram[499]  = 132;
  ram[500]  = 131;
  ram[501]  = 131;
  ram[502]  = 131;
  ram[503]  = 131;
  ram[504]  = 131;
  ram[505]  = 132;
  ram[506]  = 132;
  ram[507]  = 131;
  ram[508]  = 132;
  ram[509]  = 133;
  ram[510]  = 131;
  ram[511]  = 129;
  ram[512]  = 130;
  ram[513]  = 133;
  ram[514]  = 131;
  ram[515]  = 130;
  ram[516]  = 130;
  ram[517]  = 130;
  ram[518]  = 129;
  ram[519]  = 129;
  ram[520]  = 129;
  ram[521]  = 129;
  ram[522]  = 130;
  ram[523]  = 130;
  ram[524]  = 129;
  ram[525]  = 129;
  ram[526]  = 129;
  ram[527]  = 129;
  ram[528]  = 130;
  ram[529]  = 131;
  ram[530]  = 132;
  ram[531]  = 132;
  ram[532]  = 131;
  ram[533]  = 131;
  ram[534]  = 130;
  ram[535]  = 131;
  ram[536]  = 130;
  ram[537]  = 130;
  ram[538]  = 130;
  ram[539]  = 130;
  ram[540]  = 130;
  ram[541]  = 130;
  ram[542]  = 130;
  ram[543]  = 130;
  ram[544]  = 130;
  ram[545]  = 130;
  ram[546]  = 130;
  ram[547]  = 130;
  ram[548]  = 130;
  ram[549]  = 130;
  ram[550]  = 130;
  ram[551]  = 130;
  ram[552]  = 129;
  ram[553]  = 130;
  ram[554]  = 130;
  ram[555]  = 130;
  ram[556]  = 131;
  ram[557]  = 131;
  ram[558]  = 131;
  ram[559]  = 131;
  ram[560]  = 131;
  ram[561]  = 131;
  ram[562]  = 131;
  ram[563]  = 131;
  ram[564]  = 130;
  ram[565]  = 130;
  ram[566]  = 130;
  ram[567]  = 129;
  ram[568]  = 129;
  ram[569]  = 130;
  ram[570]  = 130;
  ram[571]  = 130;
  ram[572]  = 131;
  ram[573]  = 132;
  ram[574]  = 130;
  ram[575]  = 129;
  ram[576]  = 131;
  ram[577]  = 134;
  ram[578]  = 133;
  ram[579]  = 132;
  ram[580]  = 132;
  ram[581]  = 132;
  ram[582]  = 130;
  ram[583]  = 130;
  ram[584]  = 130;
  ram[585]  = 130;
  ram[586]  = 131;
  ram[587]  = 131;
  ram[588]  = 130;
  ram[589]  = 130;
  ram[590]  = 130;
  ram[591]  = 130;
  ram[592]  = 131;
  ram[593]  = 133;
  ram[594]  = 133;
  ram[595]  = 133;
  ram[596]  = 132;
  ram[597]  = 132;
  ram[598]  = 131;
  ram[599]  = 131;
  ram[600]  = 132;
  ram[601]  = 132;
  ram[602]  = 132;
  ram[603]  = 132;
  ram[604]  = 132;
  ram[605]  = 132;
  ram[606]  = 132;
  ram[607]  = 131;
  ram[608]  = 132;
  ram[609]  = 132;
  ram[610]  = 132;
  ram[611]  = 132;
  ram[612]  = 132;
  ram[613]  = 133;
  ram[614]  = 133;
  ram[615]  = 133;
  ram[616]  = 133;
  ram[617]  = 133;
  ram[618]  = 133;
  ram[619]  = 133;
  ram[620]  = 134;
  ram[621]  = 134;
  ram[622]  = 134;
  ram[623]  = 134;
  ram[624]  = 133;
  ram[625]  = 133;
  ram[626]  = 133;
  ram[627]  = 133;
  ram[628]  = 132;
  ram[629]  = 132;
  ram[630]  = 132;
  ram[631]  = 131;
  ram[632]  = 131;
  ram[633]  = 132;
  ram[634]  = 132;
  ram[635]  = 131;
  ram[636]  = 132;
  ram[637]  = 132;
  ram[638]  = 131;
  ram[639]  = 129;
  ram[640]  = 132;
  ram[641]  = 135;
  ram[642]  = 133;
  ram[643]  = 132;
  ram[644]  = 132;
  ram[645]  = 132;
  ram[646]  = 130;
  ram[647]  = 130;
  ram[648]  = 130;
  ram[649]  = 130;
  ram[650]  = 130;
  ram[651]  = 130;
  ram[652]  = 130;
  ram[653]  = 130;
  ram[654]  = 130;
  ram[655]  = 130;
  ram[656]  = 132;
  ram[657]  = 132;
  ram[658]  = 132;
  ram[659]  = 132;
  ram[660]  = 132;
  ram[661]  = 132;
  ram[662]  = 132;
  ram[663]  = 132;
  ram[664]  = 131;
  ram[665]  = 131;
  ram[666]  = 131;
  ram[667]  = 131;
  ram[668]  = 131;
  ram[669]  = 131;
  ram[670]  = 131;
  ram[671]  = 131;
  ram[672]  = 131;
  ram[673]  = 131;
  ram[674]  = 131;
  ram[675]  = 130;
  ram[676]  = 130;
  ram[677]  = 130;
  ram[678]  = 130;
  ram[679]  = 130;
  ram[680]  = 130;
  ram[681]  = 130;
  ram[682]  = 130;
  ram[683]  = 130;
  ram[684]  = 130;
  ram[685]  = 130;
  ram[686]  = 131;
  ram[687]  = 131;
  ram[688]  = 131;
  ram[689]  = 131;
  ram[690]  = 130;
  ram[691]  = 131;
  ram[692]  = 130;
  ram[693]  = 130;
  ram[694]  = 130;
  ram[695]  = 130;
  ram[696]  = 130;
  ram[697]  = 131;
  ram[698]  = 131;
  ram[699]  = 130;
  ram[700]  = 130;
  ram[701]  = 130;
  ram[702]  = 130;
  ram[703]  = 128;
  ram[704]  = 131;
  ram[705]  = 134;
  ram[706]  = 132;
  ram[707]  = 131;
  ram[708]  = 131;
  ram[709]  = 131;
  ram[710]  = 128;
  ram[711]  = 129;
  ram[712]  = 129;
  ram[713]  = 129;
  ram[714]  = 129;
  ram[715]  = 129;
  ram[716]  = 129;
  ram[717]  = 129;
  ram[718]  = 129;
  ram[719]  = 129;
  ram[720]  = 130;
  ram[721]  = 131;
  ram[722]  = 130;
  ram[723]  = 131;
  ram[724]  = 130;
  ram[725]  = 131;
  ram[726]  = 130;
  ram[727]  = 130;
  ram[728]  = 127;
  ram[729]  = 129;
  ram[730]  = 128;
  ram[731]  = 129;
  ram[732]  = 128;
  ram[733]  = 130;
  ram[734]  = 129;
  ram[735]  = 130;
  ram[736]  = 132;
  ram[737]  = 133;
  ram[738]  = 132;
  ram[739]  = 132;
  ram[740]  = 131;
  ram[741]  = 132;
  ram[742]  = 131;
  ram[743]  = 132;
  ram[744]  = 130;
  ram[745]  = 131;
  ram[746]  = 130;
  ram[747]  = 131;
  ram[748]  = 131;
  ram[749]  = 132;
  ram[750]  = 132;
  ram[751]  = 132;
  ram[752]  = 130;
  ram[753]  = 130;
  ram[754]  = 129;
  ram[755]  = 129;
  ram[756]  = 129;
  ram[757]  = 129;
  ram[758]  = 129;
  ram[759]  = 129;
  ram[760]  = 128;
  ram[761]  = 129;
  ram[762]  = 129;
  ram[763]  = 129;
  ram[764]  = 129;
  ram[765]  = 129;
  ram[766]  = 129;
  ram[767]  = 128;
  ram[768]  = 131;
  ram[769]  = 133;
  ram[770]  = 132;
  ram[771]  = 130;
  ram[772]  = 129;
  ram[773]  = 129;
  ram[774]  = 128;
  ram[775]  = 129;
  ram[776]  = 129;
  ram[777]  = 129;
  ram[778]  = 129;
  ram[779]  = 129;
  ram[780]  = 129;
  ram[781]  = 129;
  ram[782]  = 128;
  ram[783]  = 128;
  ram[784]  = 130;
  ram[785]  = 129;
  ram[786]  = 128;
  ram[787]  = 129;
  ram[788]  = 129;
  ram[789]  = 130;
  ram[790]  = 128;
  ram[791]  = 128;
  ram[792]  = 128;
  ram[793]  = 128;
  ram[794]  = 128;
  ram[795]  = 129;
  ram[796]  = 128;
  ram[797]  = 129;
  ram[798]  = 128;
  ram[799]  = 129;
  ram[800]  = 126;
  ram[801]  = 128;
  ram[802]  = 127;
  ram[803]  = 128;
  ram[804]  = 127;
  ram[805]  = 128;
  ram[806]  = 127;
  ram[807]  = 128;
  ram[808]  = 128;
  ram[809]  = 128;
  ram[810]  = 128;
  ram[811]  = 128;
  ram[812]  = 128;
  ram[813]  = 128;
  ram[814]  = 128;
  ram[815]  = 129;
  ram[816]  = 129;
  ram[817]  = 130;
  ram[818]  = 130;
  ram[819]  = 130;
  ram[820]  = 130;
  ram[821]  = 130;
  ram[822]  = 130;
  ram[823]  = 130;
  ram[824]  = 128;
  ram[825]  = 129;
  ram[826]  = 129;
  ram[827]  = 128;
  ram[828]  = 128;
  ram[829]  = 129;
  ram[830]  = 128;
  ram[831]  = 127;
  ram[832]  = 131;
  ram[833]  = 133;
  ram[834]  = 132;
  ram[835]  = 131;
  ram[836]  = 130;
  ram[837]  = 130;
  ram[838]  = 129;
  ram[839]  = 129;
  ram[840]  = 129;
  ram[841]  = 129;
  ram[842]  = 129;
  ram[843]  = 129;
  ram[844]  = 129;
  ram[845]  = 129;
  ram[846]  = 128;
  ram[847]  = 128;
  ram[848]  = 129;
  ram[849]  = 129;
  ram[850]  = 128;
  ram[851]  = 129;
  ram[852]  = 128;
  ram[853]  = 129;
  ram[854]  = 128;
  ram[855]  = 129;
  ram[856]  = 129;
  ram[857]  = 130;
  ram[858]  = 128;
  ram[859]  = 129;
  ram[860]  = 128;
  ram[861]  = 128;
  ram[862]  = 126;
  ram[863]  = 127;
  ram[864]  = 129;
  ram[865]  = 129;
  ram[866]  = 129;
  ram[867]  = 130;
  ram[868]  = 130;
  ram[869]  = 131;
  ram[870]  = 131;
  ram[871]  = 132;
  ram[872]  = 131;
  ram[873]  = 132;
  ram[874]  = 131;
  ram[875]  = 132;
  ram[876]  = 131;
  ram[877]  = 132;
  ram[878]  = 131;
  ram[879]  = 132;
  ram[880]  = 130;
  ram[881]  = 130;
  ram[882]  = 130;
  ram[883]  = 130;
  ram[884]  = 130;
  ram[885]  = 130;
  ram[886]  = 130;
  ram[887]  = 130;
  ram[888]  = 130;
  ram[889]  = 130;
  ram[890]  = 130;
  ram[891]  = 129;
  ram[892]  = 128;
  ram[893]  = 128;
  ram[894]  = 128;
  ram[895]  = 126;
  ram[896]  = 129;
  ram[897]  = 132;
  ram[898]  = 131;
  ram[899]  = 130;
  ram[900]  = 129;
  ram[901]  = 129;
  ram[902]  = 127;
  ram[903]  = 128;
  ram[904]  = 129;
  ram[905]  = 129;
  ram[906]  = 129;
  ram[907]  = 129;
  ram[908]  = 128;
  ram[909]  = 128;
  ram[910]  = 127;
  ram[911]  = 127;
  ram[912]  = 127;
  ram[913]  = 127;
  ram[914]  = 127;
  ram[915]  = 127;
  ram[916]  = 127;
  ram[917]  = 127;
  ram[918]  = 127;
  ram[919]  = 128;
  ram[920]  = 126;
  ram[921]  = 127;
  ram[922]  = 126;
  ram[923]  = 127;
  ram[924]  = 126;
  ram[925]  = 127;
  ram[926]  = 126;
  ram[927]  = 126;
  ram[928]  = 126;
  ram[929]  = 126;
  ram[930]  = 126;
  ram[931]  = 127;
  ram[932]  = 126;
  ram[933]  = 127;
  ram[934]  = 126;
  ram[935]  = 127;
  ram[936]  = 126;
  ram[937]  = 127;
  ram[938]  = 126;
  ram[939]  = 127;
  ram[940]  = 126;
  ram[941]  = 127;
  ram[942]  = 127;
  ram[943]  = 127;
  ram[944]  = 129;
  ram[945]  = 129;
  ram[946]  = 129;
  ram[947]  = 129;
  ram[948]  = 129;
  ram[949]  = 129;
  ram[950]  = 129;
  ram[951]  = 129;
  ram[952]  = 129;
  ram[953]  = 130;
  ram[954]  = 129;
  ram[955]  = 128;
  ram[956]  = 128;
  ram[957]  = 128;
  ram[958]  = 127;
  ram[959]  = 126;
  ram[960]  = 126;
  ram[961]  = 130;
  ram[962]  = 129;
  ram[963]  = 128;
  ram[964]  = 127;
  ram[965]  = 127;
  ram[966]  = 127;
  ram[967]  = 127;
  ram[968]  = 127;
  ram[969]  = 127;
  ram[970]  = 127;
  ram[971]  = 127;
  ram[972]  = 127;
  ram[973]  = 126;
  ram[974]  = 126;
  ram[975]  = 126;
  ram[976]  = 125;
  ram[977]  = 126;
  ram[978]  = 126;
  ram[979]  = 126;
  ram[980]  = 126;
  ram[981]  = 126;
  ram[982]  = 125;
  ram[983]  = 127;
  ram[984]  = 125;
  ram[985]  = 126;
  ram[986]  = 125;
  ram[987]  = 125;
  ram[988]  = 127;
  ram[989]  = 128;
  ram[990]  = 127;
  ram[991]  = 128;
  ram[992]  = 129;
  ram[993]  = 129;
  ram[994]  = 128;
  ram[995]  = 127;
  ram[996]  = 125;
  ram[997]  = 125;
  ram[998]  = 124;
  ram[999]  = 124;
  ram[1000]  = 126;
  ram[1001]  = 126;
  ram[1002]  = 126;
  ram[1003]  = 126;
  ram[1004]  = 126;
  ram[1005]  = 126;
  ram[1006]  = 126;
  ram[1007]  = 127;
  ram[1008]  = 127;
  ram[1009]  = 128;
  ram[1010]  = 128;
  ram[1011]  = 129;
  ram[1012]  = 129;
  ram[1013]  = 129;
  ram[1014]  = 129;
  ram[1015]  = 129;
  ram[1016]  = 126;
  ram[1017]  = 127;
  ram[1018]  = 127;
  ram[1019]  = 126;
  ram[1020]  = 126;
  ram[1021]  = 127;
  ram[1022]  = 127;
  ram[1023]  = 125;
  ram[1024]  = 127;
  ram[1025]  = 131;
  ram[1026]  = 131;
  ram[1027]  = 126;
  ram[1028]  = 127;
  ram[1029]  = 123;
  ram[1030]  = 124;
  ram[1031]  = 105;
  ram[1032]  = 111;
  ram[1033]  = 116;
  ram[1034]  = 114;
  ram[1035]  = 110;
  ram[1036]  = 113;
  ram[1037]  = 105;
  ram[1038]  = 120;
  ram[1039]  = 122;
  ram[1040]  = 116;
  ram[1041]  = 111;
  ram[1042]  = 125;
  ram[1043]  = 123;
  ram[1044]  = 128;
  ram[1045]  = 124;
  ram[1046]  = 123;
  ram[1047]  = 118;
  ram[1048]  = 110;
  ram[1049]  = 118;
  ram[1050]  = 122;
  ram[1051]  = 126;
  ram[1052]  = 125;
  ram[1053]  = 118;
  ram[1054]  = 104;
  ram[1055]  = 111;
  ram[1056]  = 113;
  ram[1057]  = 111;
  ram[1058]  = 111;
  ram[1059]  = 124;
  ram[1060]  = 125;
  ram[1061]  = 123;
  ram[1062]  = 115;
  ram[1063]  = 107;
  ram[1064]  = 115;
  ram[1065]  = 124;
  ram[1066]  = 124;
  ram[1067]  = 124;
  ram[1068]  = 120;
  ram[1069]  = 125;
  ram[1070]  = 107;
  ram[1071]  = 106;
  ram[1072]  = 124;
  ram[1073]  = 122;
  ram[1074]  = 105;
  ram[1075]  = 117;
  ram[1076]  = 106;
  ram[1077]  = 111;
  ram[1078]  = 108;
  ram[1079]  = 109;
  ram[1080]  = 109;
  ram[1081]  = 113;
  ram[1082]  = 107;
  ram[1083]  = 117;
  ram[1084]  = 127;
  ram[1085]  = 124;
  ram[1086]  = 122;
  ram[1087]  = 122;
  ram[1088]  = 124;
  ram[1089]  = 129;
  ram[1090]  = 122;
  ram[1091]  = 125;
  ram[1092]  = 130;
  ram[1093]  = 115;
  ram[1094]  = 127;
  ram[1095]  = 192;
  ram[1096]  = 176;
  ram[1097]  = 177;
  ram[1098]  = 173;
  ram[1099]  = 187;
  ram[1100]  = 168;
  ram[1101]  = 198;
  ram[1102]  = 125;
  ram[1103]  = 102;
  ram[1104]  = 183;
  ram[1105]  = 190;
  ram[1106]  = 111;
  ram[1107]  = 127;
  ram[1108]  = 122;
  ram[1109]  = 125;
  ram[1110]  = 123;
  ram[1111]  = 137;
  ram[1112]  = 195;
  ram[1113]  = 157;
  ram[1114]  = 117;
  ram[1115]  = 127;
  ram[1116]  = 112;
  ram[1117]  = 167;
  ram[1118]  = 186;
  ram[1119]  = 176;
  ram[1120]  = 179;
  ram[1121]  = 183;
  ram[1122]  = 172;
  ram[1123]  = 119;
  ram[1124]  = 122;
  ram[1125]  = 114;
  ram[1126]  = 138;
  ram[1127]  = 193;
  ram[1128]  = 148;
  ram[1129]  = 118;
  ram[1130]  = 128;
  ram[1131]  = 119;
  ram[1132]  = 127;
  ram[1133]  = 113;
  ram[1134]  = 180;
  ram[1135]  = 194;
  ram[1136]  = 104;
  ram[1137]  = 114;
  ram[1138]  = 194;
  ram[1139]  = 173;
  ram[1140]  = 181;
  ram[1141]  = 169;
  ram[1142]  = 181;
  ram[1143]  = 173;
  ram[1144]  = 180;
  ram[1145]  = 172;
  ram[1146]  = 186;
  ram[1147]  = 137;
  ram[1148]  = 119;
  ram[1149]  = 123;
  ram[1150]  = 126;
  ram[1151]  = 123;
  ram[1152]  = 128;
  ram[1153]  = 117;
  ram[1154]  = 129;
  ram[1155]  = 119;
  ram[1156]  = 114;
  ram[1157]  = 98;
  ram[1158]  = 134;
  ram[1159]  = 255;
  ram[1160]  = 250;
  ram[1161]  = 255;
  ram[1162]  = 255;
  ram[1163]  = 255;
  ram[1164]  = 255;
  ram[1165]  = 255;
  ram[1166]  = 130;
  ram[1167]  = 82;
  ram[1168]  = 255;
  ram[1169]  = 253;
  ram[1170]  = 102;
  ram[1171]  = 118;
  ram[1172]  = 122;
  ram[1173]  = 116;
  ram[1174]  = 116;
  ram[1175]  = 159;
  ram[1176]  = 255;
  ram[1177]  = 192;
  ram[1178]  = 102;
  ram[1179]  = 106;
  ram[1180]  = 96;
  ram[1181]  = 222;
  ram[1182]  = 255;
  ram[1183]  = 253;
  ram[1184]  = 254;
  ram[1185]  = 253;
  ram[1186]  = 238;
  ram[1187]  = 90;
  ram[1188]  = 100;
  ram[1189]  = 112;
  ram[1190]  = 163;
  ram[1191]  = 255;
  ram[1192]  = 171;
  ram[1193]  = 112;
  ram[1194]  = 117;
  ram[1195]  = 129;
  ram[1196]  = 99;
  ram[1197]  = 69;
  ram[1198]  = 255;
  ram[1199]  = 255;
  ram[1200]  = 76;
  ram[1201]  = 104;
  ram[1202]  = 255;
  ram[1203]  = 244;
  ram[1204]  = 255;
  ram[1205]  = 253;
  ram[1206]  = 255;
  ram[1207]  = 252;
  ram[1208]  = 254;
  ram[1209]  = 252;
  ram[1210]  = 255;
  ram[1211]  = 152;
  ram[1212]  = 117;
  ram[1213]  = 127;
  ram[1214]  = 125;
  ram[1215]  = 121;
  ram[1216]  = 117;
  ram[1217]  = 122;
  ram[1218]  = 125;
  ram[1219]  = 119;
  ram[1220]  = 124;
  ram[1221]  = 211;
  ram[1222]  = 178;
  ram[1223]  = 137;
  ram[1224]  = 137;
  ram[1225]  = 139;
  ram[1226]  = 134;
  ram[1227]  = 143;
  ram[1228]  = 141;
  ram[1229]  = 156;
  ram[1230]  = 116;
  ram[1231]  = 88;
  ram[1232]  = 240;
  ram[1233]  = 246;
  ram[1234]  = 95;
  ram[1235]  = 117;
  ram[1236]  = 122;
  ram[1237]  = 125;
  ram[1238]  = 111;
  ram[1239]  = 149;
  ram[1240]  = 255;
  ram[1241]  = 167;
  ram[1242]  = 90;
  ram[1243]  = 169;
  ram[1244]  = 213;
  ram[1245]  = 144;
  ram[1246]  = 139;
  ram[1247]  = 140;
  ram[1248]  = 140;
  ram[1249]  = 135;
  ram[1250]  = 139;
  ram[1251]  = 218;
  ram[1252]  = 183;
  ram[1253]  = 97;
  ram[1254]  = 150;
  ram[1255]  = 252;
  ram[1256]  = 163;
  ram[1257]  = 111;
  ram[1258]  = 118;
  ram[1259]  = 104;
  ram[1260]  = 191;
  ram[1261]  = 215;
  ram[1262]  = 130;
  ram[1263]  = 143;
  ram[1264]  = 100;
  ram[1265]  = 106;
  ram[1266]  = 254;
  ram[1267]  = 207;
  ram[1268]  = 127;
  ram[1269]  = 137;
  ram[1270]  = 150;
  ram[1271]  = 138;
  ram[1272]  = 144;
  ram[1273]  = 142;
  ram[1274]  = 149;
  ram[1275]  = 120;
  ram[1276]  = 124;
  ram[1277]  = 124;
  ram[1278]  = 118;
  ram[1279]  = 123;
  ram[1280]  = 120;
  ram[1281]  = 125;
  ram[1282]  = 120;
  ram[1283]  = 118;
  ram[1284]  = 129;
  ram[1285]  = 250;
  ram[1286]  = 226;
  ram[1287]  = 80;
  ram[1288]  = 103;
  ram[1289]  = 105;
  ram[1290]  = 107;
  ram[1291]  = 101;
  ram[1292]  = 112;
  ram[1293]  = 111;
  ram[1294]  = 115;
  ram[1295]  = 87;
  ram[1296]  = 248;
  ram[1297]  = 251;
  ram[1298]  = 70;
  ram[1299]  = 96;
  ram[1300]  = 126;
  ram[1301]  = 122;
  ram[1302]  = 119;
  ram[1303]  = 148;
  ram[1304]  = 252;
  ram[1305]  = 184;
  ram[1306]  = 84;
  ram[1307]  = 194;
  ram[1308]  = 255;
  ram[1309]  = 134;
  ram[1310]  = 91;
  ram[1311]  = 100;
  ram[1312]  = 107;
  ram[1313]  = 99;
  ram[1314]  = 119;
  ram[1315]  = 244;
  ram[1316]  = 211;
  ram[1317]  = 90;
  ram[1318]  = 162;
  ram[1319]  = 255;
  ram[1320]  = 162;
  ram[1321]  = 108;
  ram[1322]  = 98;
  ram[1323]  = 65;
  ram[1324]  = 250;
  ram[1325]  = 255;
  ram[1326]  = 92;
  ram[1327]  = 105;
  ram[1328]  = 111;
  ram[1329]  = 108;
  ram[1330]  = 255;
  ram[1331]  = 218;
  ram[1332]  = 80;
  ram[1333]  = 103;
  ram[1334]  = 105;
  ram[1335]  = 106;
  ram[1336]  = 108;
  ram[1337]  = 110;
  ram[1338]  = 112;
  ram[1339]  = 116;
  ram[1340]  = 121;
  ram[1341]  = 121;
  ram[1342]  = 125;
  ram[1343]  = 121;
  ram[1344]  = 119;
  ram[1345]  = 125;
  ram[1346]  = 120;
  ram[1347]  = 121;
  ram[1348]  = 118;
  ram[1349]  = 251;
  ram[1350]  = 198;
  ram[1351]  = 106;
  ram[1352]  = 115;
  ram[1353]  = 116;
  ram[1354]  = 120;
  ram[1355]  = 116;
  ram[1356]  = 111;
  ram[1357]  = 126;
  ram[1358]  = 120;
  ram[1359]  = 86;
  ram[1360]  = 236;
  ram[1361]  = 228;
  ram[1362]  = 214;
  ram[1363]  = 227;
  ram[1364]  = 99;
  ram[1365]  = 117;
  ram[1366]  = 109;
  ram[1367]  = 151;
  ram[1368]  = 253;
  ram[1369]  = 163;
  ram[1370]  = 85;
  ram[1371]  = 183;
  ram[1372]  = 242;
  ram[1373]  = 135;
  ram[1374]  = 107;
  ram[1375]  = 113;
  ram[1376]  = 115;
  ram[1377]  = 117;
  ram[1378]  = 126;
  ram[1379]  = 236;
  ram[1380]  = 196;
  ram[1381]  = 84;
  ram[1382]  = 152;
  ram[1383]  = 254;
  ram[1384]  = 153;
  ram[1385]  = 89;
  ram[1386]  = 189;
  ram[1387]  = 238;
  ram[1388]  = 118;
  ram[1389]  = 117;
  ram[1390]  = 108;
  ram[1391]  = 112;
  ram[1392]  = 118;
  ram[1393]  = 92;
  ram[1394]  = 252;
  ram[1395]  = 214;
  ram[1396]  = 85;
  ram[1397]  = 121;
  ram[1398]  = 118;
  ram[1399]  = 115;
  ram[1400]  = 113;
  ram[1401]  = 116;
  ram[1402]  = 118;
  ram[1403]  = 119;
  ram[1404]  = 125;
  ram[1405]  = 116;
  ram[1406]  = 118;
  ram[1407]  = 115;
  ram[1408]  = 119;
  ram[1409]  = 123;
  ram[1410]  = 119;
  ram[1411]  = 120;
  ram[1412]  = 124;
  ram[1413]  = 251;
  ram[1414]  = 200;
  ram[1415]  = 60;
  ram[1416]  = 92;
  ram[1417]  = 93;
  ram[1418]  = 88;
  ram[1419]  = 93;
  ram[1420]  = 107;
  ram[1421]  = 119;
  ram[1422]  = 120;
  ram[1423]  = 89;
  ram[1424]  = 241;
  ram[1425]  = 236;
  ram[1426]  = 255;
  ram[1427]  = 255;
  ram[1428]  = 63;
  ram[1429]  = 100;
  ram[1430]  = 100;
  ram[1431]  = 149;
  ram[1432]  = 254;
  ram[1433]  = 174;
  ram[1434]  = 83;
  ram[1435]  = 193;
  ram[1436]  = 251;
  ram[1437]  = 113;
  ram[1438]  = 71;
  ram[1439]  = 81;
  ram[1440]  = 88;
  ram[1441]  = 75;
  ram[1442]  = 108;
  ram[1443]  = 242;
  ram[1444]  = 203;
  ram[1445]  = 82;
  ram[1446]  = 153;
  ram[1447]  = 255;
  ram[1448]  = 140;
  ram[1449]  = 32;
  ram[1450]  = 213;
  ram[1451]  = 255;
  ram[1452]  = 109;
  ram[1453]  = 101;
  ram[1454]  = 113;
  ram[1455]  = 124;
  ram[1456]  = 113;
  ram[1457]  = 109;
  ram[1458]  = 255;
  ram[1459]  = 207;
  ram[1460]  = 51;
  ram[1461]  = 90;
  ram[1462]  = 88;
  ram[1463]  = 87;
  ram[1464]  = 89;
  ram[1465]  = 102;
  ram[1466]  = 115;
  ram[1467]  = 116;
  ram[1468]  = 120;
  ram[1469]  = 119;
  ram[1470]  = 123;
  ram[1471]  = 120;
  ram[1472]  = 118;
  ram[1473]  = 117;
  ram[1474]  = 123;
  ram[1475]  = 113;
  ram[1476]  = 120;
  ram[1477]  = 236;
  ram[1478]  = 221;
  ram[1479]  = 245;
  ram[1480]  = 233;
  ram[1481]  = 249;
  ram[1482]  = 239;
  ram[1483]  = 255;
  ram[1484]  = 148;
  ram[1485]  = 108;
  ram[1486]  = 115;
  ram[1487]  = 80;
  ram[1488]  = 241;
  ram[1489]  = 246;
  ram[1490]  = 59;
  ram[1491]  = 80;
  ram[1492]  = 255;
  ram[1493]  = 225;
  ram[1494]  = 84;
  ram[1495]  = 138;
  ram[1496]  = 253;
  ram[1497]  = 166;
  ram[1498]  = 72;
  ram[1499]  = 184;
  ram[1500]  = 237;
  ram[1501]  = 231;
  ram[1502]  = 249;
  ram[1503]  = 241;
  ram[1504]  = 241;
  ram[1505]  = 248;
  ram[1506]  = 227;
  ram[1507]  = 232;
  ram[1508]  = 193;
  ram[1509]  = 76;
  ram[1510]  = 152;
  ram[1511]  = 235;
  ram[1512]  = 212;
  ram[1513]  = 255;
  ram[1514]  = 111;
  ram[1515]  = 83;
  ram[1516]  = 98;
  ram[1517]  = 112;
  ram[1518]  = 118;
  ram[1519]  = 110;
  ram[1520]  = 114;
  ram[1521]  = 102;
  ram[1522]  = 250;
  ram[1523]  = 219;
  ram[1524]  = 244;
  ram[1525]  = 233;
  ram[1526]  = 242;
  ram[1527]  = 239;
  ram[1528]  = 249;
  ram[1529]  = 160;
  ram[1530]  = 105;
  ram[1531]  = 117;
  ram[1532]  = 119;
  ram[1533]  = 115;
  ram[1534]  = 118;
  ram[1535]  = 112;
  ram[1536]  = 116;
  ram[1537]  = 120;
  ram[1538]  = 118;
  ram[1539]  = 115;
  ram[1540]  = 124;
  ram[1541]  = 248;
  ram[1542]  = 248;
  ram[1543]  = 250;
  ram[1544]  = 249;
  ram[1545]  = 251;
  ram[1546]  = 246;
  ram[1547]  = 255;
  ram[1548]  = 125;
  ram[1549]  = 73;
  ram[1550]  = 106;
  ram[1551]  = 76;
  ram[1552]  = 244;
  ram[1553]  = 249;
  ram[1554]  = 69;
  ram[1555]  = 102;
  ram[1556]  = 255;
  ram[1557]  = 220;
  ram[1558]  = 49;
  ram[1559]  = 120;
  ram[1560]  = 244;
  ram[1561]  = 174;
  ram[1562]  = 78;
  ram[1563]  = 184;
  ram[1564]  = 236;
  ram[1565]  = 247;
  ram[1566]  = 249;
  ram[1567]  = 255;
  ram[1568]  = 255;
  ram[1569]  = 254;
  ram[1570]  = 244;
  ram[1571]  = 236;
  ram[1572]  = 197;
  ram[1573]  = 83;
  ram[1574]  = 147;
  ram[1575]  = 237;
  ram[1576]  = 231;
  ram[1577]  = 255;
  ram[1578]  = 110;
  ram[1579]  = 66;
  ram[1580]  = 102;
  ram[1581]  = 111;
  ram[1582]  = 109;
  ram[1583]  = 116;
  ram[1584]  = 110;
  ram[1585]  = 102;
  ram[1586]  = 250;
  ram[1587]  = 228;
  ram[1588]  = 255;
  ram[1589]  = 250;
  ram[1590]  = 255;
  ram[1591]  = 250;
  ram[1592]  = 252;
  ram[1593]  = 151;
  ram[1594]  = 106;
  ram[1595]  = 113;
  ram[1596]  = 121;
  ram[1597]  = 121;
  ram[1598]  = 113;
  ram[1599]  = 114;
  ram[1600]  = 117;
  ram[1601]  = 112;
  ram[1602]  = 114;
  ram[1603]  = 112;
  ram[1604]  = 114;
  ram[1605]  = 84;
  ram[1606]  = 75;
  ram[1607]  = 81;
  ram[1608]  = 69;
  ram[1609]  = 78;
  ram[1610]  = 70;
  ram[1611]  = 48;
  ram[1612]  = 189;
  ram[1613]  = 255;
  ram[1614]  = 121;
  ram[1615]  = 63;
  ram[1616]  = 239;
  ram[1617]  = 251;
  ram[1618]  = 81;
  ram[1619]  = 100;
  ram[1620]  = 67;
  ram[1621]  = 101;
  ram[1622]  = 255;
  ram[1623]  = 236;
  ram[1624]  = 230;
  ram[1625]  = 166;
  ram[1626]  = 66;
  ram[1627]  = 181;
  ram[1628]  = 242;
  ram[1629]  = 109;
  ram[1630]  = 73;
  ram[1631]  = 74;
  ram[1632]  = 76;
  ram[1633]  = 79;
  ram[1634]  = 96;
  ram[1635]  = 237;
  ram[1636]  = 199;
  ram[1637]  = 81;
  ram[1638]  = 147;
  ram[1639]  = 255;
  ram[1640]  = 131;
  ram[1641]  = 41;
  ram[1642]  = 200;
  ram[1643]  = 255;
  ram[1644]  = 125;
  ram[1645]  = 96;
  ram[1646]  = 112;
  ram[1647]  = 111;
  ram[1648]  = 112;
  ram[1649]  = 97;
  ram[1650]  = 255;
  ram[1651]  = 198;
  ram[1652]  = 48;
  ram[1653]  = 77;
  ram[1654]  = 78;
  ram[1655]  = 78;
  ram[1656]  = 83;
  ram[1657]  = 101;
  ram[1658]  = 110;
  ram[1659]  = 113;
  ram[1660]  = 115;
  ram[1661]  = 112;
  ram[1662]  = 115;
  ram[1663]  = 110;
  ram[1664]  = 112;
  ram[1665]  = 114;
  ram[1666]  = 118;
  ram[1667]  = 115;
  ram[1668]  = 103;
  ram[1669]  = 110;
  ram[1670]  = 107;
  ram[1671]  = 106;
  ram[1672]  = 108;
  ram[1673]  = 106;
  ram[1674]  = 105;
  ram[1675]  = 85;
  ram[1676]  = 189;
  ram[1677]  = 255;
  ram[1678]  = 108;
  ram[1679]  = 66;
  ram[1680]  = 242;
  ram[1681]  = 245;
  ram[1682]  = 85;
  ram[1683]  = 103;
  ram[1684]  = 96;
  ram[1685]  = 128;
  ram[1686]  = 250;
  ram[1687]  = 228;
  ram[1688]  = 235;
  ram[1689]  = 163;
  ram[1690]  = 72;
  ram[1691]  = 186;
  ram[1692]  = 248;
  ram[1693]  = 127;
  ram[1694]  = 101;
  ram[1695]  = 102;
  ram[1696]  = 107;
  ram[1697]  = 102;
  ram[1698]  = 110;
  ram[1699]  = 249;
  ram[1700]  = 196;
  ram[1701]  = 72;
  ram[1702]  = 150;
  ram[1703]  = 254;
  ram[1704]  = 150;
  ram[1705]  = 62;
  ram[1706]  = 202;
  ram[1707]  = 250;
  ram[1708]  = 105;
  ram[1709]  = 99;
  ram[1710]  = 113;
  ram[1711]  = 112;
  ram[1712]  = 105;
  ram[1713]  = 100;
  ram[1714]  = 251;
  ram[1715]  = 212;
  ram[1716]  = 78;
  ram[1717]  = 104;
  ram[1718]  = 104;
  ram[1719]  = 108;
  ram[1720]  = 104;
  ram[1721]  = 109;
  ram[1722]  = 108;
  ram[1723]  = 113;
  ram[1724]  = 113;
  ram[1725]  = 114;
  ram[1726]  = 112;
  ram[1727]  = 112;
  ram[1728]  = 110;
  ram[1729]  = 117;
  ram[1730]  = 107;
  ram[1731]  = 112;
  ram[1732]  = 115;
  ram[1733]  = 110;
  ram[1734]  = 109;
  ram[1735]  = 105;
  ram[1736]  = 105;
  ram[1737]  = 95;
  ram[1738]  = 103;
  ram[1739]  = 75;
  ram[1740]  = 189;
  ram[1741]  = 253;
  ram[1742]  = 109;
  ram[1743]  = 59;
  ram[1744]  = 247;
  ram[1745]  = 253;
  ram[1746]  = 82;
  ram[1747]  = 105;
  ram[1748]  = 115;
  ram[1749]  = 101;
  ram[1750]  = 62;
  ram[1751]  = 119;
  ram[1752]  = 254;
  ram[1753]  = 170;
  ram[1754]  = 73;
  ram[1755]  = 181;
  ram[1756]  = 252;
  ram[1757]  = 128;
  ram[1758]  = 102;
  ram[1759]  = 104;
  ram[1760]  = 112;
  ram[1761]  = 101;
  ram[1762]  = 124;
  ram[1763]  = 236;
  ram[1764]  = 206;
  ram[1765]  = 75;
  ram[1766]  = 149;
  ram[1767]  = 255;
  ram[1768]  = 156;
  ram[1769]  = 91;
  ram[1770]  = 81;
  ram[1771]  = 43;
  ram[1772]  = 234;
  ram[1773]  = 255;
  ram[1774]  = 94;
  ram[1775]  = 100;
  ram[1776]  = 110;
  ram[1777]  = 91;
  ram[1778]  = 252;
  ram[1779]  = 212;
  ram[1780]  = 65;
  ram[1781]  = 105;
  ram[1782]  = 108;
  ram[1783]  = 104;
  ram[1784]  = 107;
  ram[1785]  = 104;
  ram[1786]  = 103;
  ram[1787]  = 111;
  ram[1788]  = 110;
  ram[1789]  = 112;
  ram[1790]  = 108;
  ram[1791]  = 108;
  ram[1792]  = 111;
  ram[1793]  = 106;
  ram[1794]  = 117;
  ram[1795]  = 108;
  ram[1796]  = 107;
  ram[1797]  = 122;
  ram[1798]  = 118;
  ram[1799]  = 128;
  ram[1800]  = 120;
  ram[1801]  = 118;
  ram[1802]  = 119;
  ram[1803]  = 106;
  ram[1804]  = 179;
  ram[1805]  = 243;
  ram[1806]  = 101;
  ram[1807]  = 62;
  ram[1808]  = 238;
  ram[1809]  = 248;
  ram[1810]  = 82;
  ram[1811]  = 107;
  ram[1812]  = 99;
  ram[1813]  = 113;
  ram[1814]  = 98;
  ram[1815]  = 138;
  ram[1816]  = 254;
  ram[1817]  = 162;
  ram[1818]  = 75;
  ram[1819]  = 183;
  ram[1820]  = 244;
  ram[1821]  = 132;
  ram[1822]  = 95;
  ram[1823]  = 107;
  ram[1824]  = 101;
  ram[1825]  = 107;
  ram[1826]  = 114;
  ram[1827]  = 241;
  ram[1828]  = 195;
  ram[1829]  = 81;
  ram[1830]  = 140;
  ram[1831]  = 255;
  ram[1832]  = 151;
  ram[1833]  = 93;
  ram[1834]  = 99;
  ram[1835]  = 82;
  ram[1836]  = 210;
  ram[1837]  = 231;
  ram[1838]  = 96;
  ram[1839]  = 124;
  ram[1840]  = 95;
  ram[1841]  = 85;
  ram[1842]  = 254;
  ram[1843]  = 199;
  ram[1844]  = 98;
  ram[1845]  = 115;
  ram[1846]  = 123;
  ram[1847]  = 117;
  ram[1848]  = 121;
  ram[1849]  = 124;
  ram[1850]  = 127;
  ram[1851]  = 107;
  ram[1852]  = 111;
  ram[1853]  = 107;
  ram[1854]  = 108;
  ram[1855]  = 109;
  ram[1856]  = 108;
  ram[1857]  = 107;
  ram[1858]  = 103;
  ram[1859]  = 107;
  ram[1860]  = 118;
  ram[1861]  = 255;
  ram[1862]  = 255;
  ram[1863]  = 253;
  ram[1864]  = 250;
  ram[1865]  = 255;
  ram[1866]  = 247;
  ram[1867]  = 255;
  ram[1868]  = 114;
  ram[1869]  = 59;
  ram[1870]  = 100;
  ram[1871]  = 63;
  ram[1872]  = 255;
  ram[1873]  = 251;
  ram[1874]  = 82;
  ram[1875]  = 108;
  ram[1876]  = 110;
  ram[1877]  = 104;
  ram[1878]  = 99;
  ram[1879]  = 144;
  ram[1880]  = 252;
  ram[1881]  = 177;
  ram[1882]  = 67;
  ram[1883]  = 193;
  ram[1884]  = 255;
  ram[1885]  = 136;
  ram[1886]  = 101;
  ram[1887]  = 108;
  ram[1888]  = 100;
  ram[1889]  = 106;
  ram[1890]  = 129;
  ram[1891]  = 250;
  ram[1892]  = 206;
  ram[1893]  = 70;
  ram[1894]  = 151;
  ram[1895]  = 255;
  ram[1896]  = 154;
  ram[1897]  = 90;
  ram[1898]  = 106;
  ram[1899]  = 107;
  ram[1900]  = 82;
  ram[1901]  = 35;
  ram[1902]  = 255;
  ram[1903]  = 255;
  ram[1904]  = 52;
  ram[1905]  = 95;
  ram[1906]  = 255;
  ram[1907]  = 233;
  ram[1908]  = 253;
  ram[1909]  = 255;
  ram[1910]  = 251;
  ram[1911]  = 255;
  ram[1912]  = 253;
  ram[1913]  = 253;
  ram[1914]  = 255;
  ram[1915]  = 140;
  ram[1916]  = 100;
  ram[1917]  = 105;
  ram[1918]  = 108;
  ram[1919]  = 103;
  ram[1920]  = 103;
  ram[1921]  = 106;
  ram[1922]  = 109;
  ram[1923]  = 100;
  ram[1924]  = 107;
  ram[1925]  = 201;
  ram[1926]  = 172;
  ram[1927]  = 194;
  ram[1928]  = 179;
  ram[1929]  = 197;
  ram[1930]  = 178;
  ram[1931]  = 205;
  ram[1932]  = 118;
  ram[1933]  = 93;
  ram[1934]  = 93;
  ram[1935]  = 84;
  ram[1936]  = 194;
  ram[1937]  = 206;
  ram[1938]  = 88;
  ram[1939]  = 101;
  ram[1940]  = 102;
  ram[1941]  = 109;
  ram[1942]  = 97;
  ram[1943]  = 125;
  ram[1944]  = 219;
  ram[1945]  = 133;
  ram[1946]  = 80;
  ram[1947]  = 158;
  ram[1948]  = 206;
  ram[1949]  = 116;
  ram[1950]  = 98;
  ram[1951]  = 99;
  ram[1952]  = 107;
  ram[1953]  = 100;
  ram[1954]  = 110;
  ram[1955]  = 207;
  ram[1956]  = 166;
  ram[1957]  = 83;
  ram[1958]  = 127;
  ram[1959]  = 211;
  ram[1960]  = 131;
  ram[1961]  = 92;
  ram[1962]  = 98;
  ram[1963]  = 106;
  ram[1964]  = 104;
  ram[1965]  = 81;
  ram[1966]  = 198;
  ram[1967]  = 215;
  ram[1968]  = 70;
  ram[1969]  = 91;
  ram[1970]  = 217;
  ram[1971]  = 176;
  ram[1972]  = 195;
  ram[1973]  = 182;
  ram[1974]  = 196;
  ram[1975]  = 182;
  ram[1976]  = 195;
  ram[1977]  = 178;
  ram[1978]  = 197;
  ram[1979]  = 124;
  ram[1980]  = 101;
  ram[1981]  = 107;
  ram[1982]  = 102;
  ram[1983]  = 104;
  ram[1984]  = 102;
  ram[1985]  = 103;
  ram[1986]  = 104;
  ram[1987]  = 106;
  ram[1988]  = 99;
  ram[1989]  = 80;
  ram[1990]  = 77;
  ram[1991]  = 73;
  ram[1992]  = 72;
  ram[1993]  = 72;
  ram[1994]  = 75;
  ram[1995]  = 76;
  ram[1996]  = 89;
  ram[1997]  = 101;
  ram[1998]  = 105;
  ram[1999]  = 98;
  ram[2000]  = 81;
  ram[2001]  = 76;
  ram[2002]  = 105;
  ram[2003]  = 103;
  ram[2004]  = 106;
  ram[2005]  = 103;
  ram[2006]  = 104;
  ram[2007]  = 87;
  ram[2008]  = 70;
  ram[2009]  = 92;
  ram[2010]  = 100;
  ram[2011]  = 81;
  ram[2012]  = 82;
  ram[2013]  = 97;
  ram[2014]  = 101;
  ram[2015]  = 103;
  ram[2016]  = 101;
  ram[2017]  = 103;
  ram[2018]  = 101;
  ram[2019]  = 76;
  ram[2020]  = 84;
  ram[2021]  = 99;
  ram[2022]  = 91;
  ram[2023]  = 76;
  ram[2024]  = 89;
  ram[2025]  = 100;
  ram[2026]  = 104;
  ram[2027]  = 106;
  ram[2028]  = 103;
  ram[2029]  = 101;
  ram[2030]  = 78;
  ram[2031]  = 74;
  ram[2032]  = 102;
  ram[2033]  = 96;
  ram[2034]  = 75;
  ram[2035]  = 83;
  ram[2036]  = 74;
  ram[2037]  = 72;
  ram[2038]  = 76;
  ram[2039]  = 78;
  ram[2040]  = 76;
  ram[2041]  = 77;
  ram[2042]  = 76;
  ram[2043]  = 88;
  ram[2044]  = 107;
  ram[2045]  = 103;
  ram[2046]  = 101;
  ram[2047]  = 100;
  ram[2048]  = 102;
  ram[2049]  = 102;
  ram[2050]  = 101;
  ram[2051]  = 100;
  ram[2052]  = 99;
  ram[2053]  = 99;
  ram[2054]  = 100;
  ram[2055]  = 100;
  ram[2056]  = 100;
  ram[2057]  = 102;
  ram[2058]  = 103;
  ram[2059]  = 102;
  ram[2060]  = 101;
  ram[2061]  = 101;
  ram[2062]  = 100;
  ram[2063]  = 99;
  ram[2064]  = 98;
  ram[2065]  = 99;
  ram[2066]  = 101;
  ram[2067]  = 102;
  ram[2068]  = 102;
  ram[2069]  = 101;
  ram[2070]  = 101;
  ram[2071]  = 101;
  ram[2072]  = 101;
  ram[2073]  = 101;
  ram[2074]  = 101;
  ram[2075]  = 102;
  ram[2076]  = 102;
  ram[2077]  = 102;
  ram[2078]  = 101;
  ram[2079]  = 101;
  ram[2080]  = 102;
  ram[2081]  = 102;
  ram[2082]  = 103;
  ram[2083]  = 105;
  ram[2084]  = 103;
  ram[2085]  = 101;
  ram[2086]  = 100;
  ram[2087]  = 100;
  ram[2088]  = 100;
  ram[2089]  = 101;
  ram[2090]  = 102;
  ram[2091]  = 103;
  ram[2092]  = 100;
  ram[2093]  = 100;
  ram[2094]  = 98;
  ram[2095]  = 98;
  ram[2096]  = 92;
  ram[2097]  = 96;
  ram[2098]  = 99;
  ram[2099]  = 102;
  ram[2100]  = 100;
  ram[2101]  = 101;
  ram[2102]  = 101;
  ram[2103]  = 102;
  ram[2104]  = 103;
  ram[2105]  = 103;
  ram[2106]  = 103;
  ram[2107]  = 103;
  ram[2108]  = 102;
  ram[2109]  = 101;
  ram[2110]  = 100;
  ram[2111]  = 100;
  ram[2112]  = 100;
  ram[2113]  = 100;
  ram[2114]  = 98;
  ram[2115]  = 98;
  ram[2116]  = 98;
  ram[2117]  = 98;
  ram[2118]  = 98;
  ram[2119]  = 100;
  ram[2120]  = 99;
  ram[2121]  = 100;
  ram[2122]  = 100;
  ram[2123]  = 98;
  ram[2124]  = 98;
  ram[2125]  = 99;
  ram[2126]  = 100;
  ram[2127]  = 98;
  ram[2128]  = 98;
  ram[2129]  = 99;
  ram[2130]  = 99;
  ram[2131]  = 100;
  ram[2132]  = 101;
  ram[2133]  = 101;
  ram[2134]  = 100;
  ram[2135]  = 100;
  ram[2136]  = 99;
  ram[2137]  = 99;
  ram[2138]  = 99;
  ram[2139]  = 99;
  ram[2140]  = 99;
  ram[2141]  = 99;
  ram[2142]  = 99;
  ram[2143]  = 99;
  ram[2144]  = 99;
  ram[2145]  = 98;
  ram[2146]  = 99;
  ram[2147]  = 100;
  ram[2148]  = 99;
  ram[2149]  = 98;
  ram[2150]  = 98;
  ram[2151]  = 99;
  ram[2152]  = 99;
  ram[2153]  = 99;
  ram[2154]  = 100;
  ram[2155]  = 100;
  ram[2156]  = 100;
  ram[2157]  = 99;
  ram[2158]  = 98;
  ram[2159]  = 98;
  ram[2160]  = 96;
  ram[2161]  = 97;
  ram[2162]  = 98;
  ram[2163]  = 98;
  ram[2164]  = 98;
  ram[2165]  = 99;
  ram[2166]  = 99;
  ram[2167]  = 99;
  ram[2168]  = 99;
  ram[2169]  = 100;
  ram[2170]  = 100;
  ram[2171]  = 100;
  ram[2172]  = 99;
  ram[2173]  = 99;
  ram[2174]  = 97;
  ram[2175]  = 98;
  ram[2176]  = 99;
  ram[2177]  = 99;
  ram[2178]  = 98;
  ram[2179]  = 98;
  ram[2180]  = 98;
  ram[2181]  = 98;
  ram[2182]  = 97;
  ram[2183]  = 98;
  ram[2184]  = 99;
  ram[2185]  = 99;
  ram[2186]  = 98;
  ram[2187]  = 97;
  ram[2188]  = 96;
  ram[2189]  = 98;
  ram[2190]  = 99;
  ram[2191]  = 98;
  ram[2192]  = 95;
  ram[2193]  = 96;
  ram[2194]  = 96;
  ram[2195]  = 96;
  ram[2196]  = 97;
  ram[2197]  = 97;
  ram[2198]  = 96;
  ram[2199]  = 96;
  ram[2200]  = 97;
  ram[2201]  = 97;
  ram[2202]  = 96;
  ram[2203]  = 96;
  ram[2204]  = 97;
  ram[2205]  = 97;
  ram[2206]  = 97;
  ram[2207]  = 97;
  ram[2208]  = 98;
  ram[2209]  = 97;
  ram[2210]  = 97;
  ram[2211]  = 97;
  ram[2212]  = 98;
  ram[2213]  = 97;
  ram[2214]  = 98;
  ram[2215]  = 98;
  ram[2216]  = 98;
  ram[2217]  = 98;
  ram[2218]  = 99;
  ram[2219]  = 99;
  ram[2220]  = 100;
  ram[2221]  = 100;
  ram[2222]  = 98;
  ram[2223]  = 99;
  ram[2224]  = 101;
  ram[2225]  = 99;
  ram[2226]  = 97;
  ram[2227]  = 97;
  ram[2228]  = 98;
  ram[2229]  = 98;
  ram[2230]  = 98;
  ram[2231]  = 97;
  ram[2232]  = 97;
  ram[2233]  = 99;
  ram[2234]  = 99;
  ram[2235]  = 99;
  ram[2236]  = 98;
  ram[2237]  = 97;
  ram[2238]  = 96;
  ram[2239]  = 96;
  ram[2240]  = 98;
  ram[2241]  = 98;
  ram[2242]  = 98;
  ram[2243]  = 98;
  ram[2244]  = 97;
  ram[2245]  = 97;
  ram[2246]  = 95;
  ram[2247]  = 95;
  ram[2248]  = 97;
  ram[2249]  = 97;
  ram[2250]  = 95;
  ram[2251]  = 95;
  ram[2252]  = 94;
  ram[2253]  = 96;
  ram[2254]  = 97;
  ram[2255]  = 96;
  ram[2256]  = 93;
  ram[2257]  = 93;
  ram[2258]  = 93;
  ram[2259]  = 94;
  ram[2260]  = 93;
  ram[2261]  = 94;
  ram[2262]  = 94;
  ram[2263]  = 94;
  ram[2264]  = 95;
  ram[2265]  = 96;
  ram[2266]  = 95;
  ram[2267]  = 96;
  ram[2268]  = 96;
  ram[2269]  = 96;
  ram[2270]  = 97;
  ram[2271]  = 97;
  ram[2272]  = 97;
  ram[2273]  = 96;
  ram[2274]  = 96;
  ram[2275]  = 96;
  ram[2276]  = 97;
  ram[2277]  = 96;
  ram[2278]  = 97;
  ram[2279]  = 98;
  ram[2280]  = 97;
  ram[2281]  = 97;
  ram[2282]  = 97;
  ram[2283]  = 98;
  ram[2284]  = 98;
  ram[2285]  = 98;
  ram[2286]  = 97;
  ram[2287]  = 95;
  ram[2288]  = 98;
  ram[2289]  = 97;
  ram[2290]  = 95;
  ram[2291]  = 95;
  ram[2292]  = 96;
  ram[2293]  = 97;
  ram[2294]  = 96;
  ram[2295]  = 96;
  ram[2296]  = 94;
  ram[2297]  = 96;
  ram[2298]  = 96;
  ram[2299]  = 97;
  ram[2300]  = 95;
  ram[2301]  = 95;
  ram[2302]  = 94;
  ram[2303]  = 94;
  ram[2304]  = 95;
  ram[2305]  = 95;
  ram[2306]  = 95;
  ram[2307]  = 95;
  ram[2308]  = 95;
  ram[2309]  = 94;
  ram[2310]  = 94;
  ram[2311]  = 93;
  ram[2312]  = 94;
  ram[2313]  = 94;
  ram[2314]  = 94;
  ram[2315]  = 94;
  ram[2316]  = 94;
  ram[2317]  = 93;
  ram[2318]  = 94;
  ram[2319]  = 94;
  ram[2320]  = 94;
  ram[2321]  = 94;
  ram[2322]  = 94;
  ram[2323]  = 94;
  ram[2324]  = 93;
  ram[2325]  = 94;
  ram[2326]  = 94;
  ram[2327]  = 93;
  ram[2328]  = 94;
  ram[2329]  = 94;
  ram[2330]  = 93;
  ram[2331]  = 94;
  ram[2332]  = 94;
  ram[2333]  = 94;
  ram[2334]  = 95;
  ram[2335]  = 95;
  ram[2336]  = 96;
  ram[2337]  = 95;
  ram[2338]  = 94;
  ram[2339]  = 94;
  ram[2340]  = 95;
  ram[2341]  = 95;
  ram[2342]  = 95;
  ram[2343]  = 97;
  ram[2344]  = 94;
  ram[2345]  = 94;
  ram[2346]  = 94;
  ram[2347]  = 95;
  ram[2348]  = 96;
  ram[2349]  = 96;
  ram[2350]  = 93;
  ram[2351]  = 93;
  ram[2352]  = 94;
  ram[2353]  = 93;
  ram[2354]  = 93;
  ram[2355]  = 93;
  ram[2356]  = 93;
  ram[2357]  = 93;
  ram[2358]  = 93;
  ram[2359]  = 93;
  ram[2360]  = 93;
  ram[2361]  = 93;
  ram[2362]  = 94;
  ram[2363]  = 94;
  ram[2364]  = 94;
  ram[2365]  = 93;
  ram[2366]  = 92;
  ram[2367]  = 91;
  ram[2368]  = 93;
  ram[2369]  = 93;
  ram[2370]  = 94;
  ram[2371]  = 94;
  ram[2372]  = 95;
  ram[2373]  = 94;
  ram[2374]  = 94;
  ram[2375]  = 93;
  ram[2376]  = 93;
  ram[2377]  = 93;
  ram[2378]  = 93;
  ram[2379]  = 94;
  ram[2380]  = 94;
  ram[2381]  = 93;
  ram[2382]  = 93;
  ram[2383]  = 93;
  ram[2384]  = 93;
  ram[2385]  = 93;
  ram[2386]  = 93;
  ram[2387]  = 93;
  ram[2388]  = 93;
  ram[2389]  = 94;
  ram[2390]  = 94;
  ram[2391]  = 93;
  ram[2392]  = 91;
  ram[2393]  = 92;
  ram[2394]  = 91;
  ram[2395]  = 92;
  ram[2396]  = 92;
  ram[2397]  = 93;
  ram[2398]  = 94;
  ram[2399]  = 94;
  ram[2400]  = 94;
  ram[2401]  = 93;
  ram[2402]  = 92;
  ram[2403]  = 93;
  ram[2404]  = 94;
  ram[2405]  = 93;
  ram[2406]  = 93;
  ram[2407]  = 94;
  ram[2408]  = 93;
  ram[2409]  = 93;
  ram[2410]  = 92;
  ram[2411]  = 94;
  ram[2412]  = 95;
  ram[2413]  = 95;
  ram[2414]  = 93;
  ram[2415]  = 93;
  ram[2416]  = 91;
  ram[2417]  = 93;
  ram[2418]  = 94;
  ram[2419]  = 94;
  ram[2420]  = 94;
  ram[2421]  = 93;
  ram[2422]  = 93;
  ram[2423]  = 93;
  ram[2424]  = 93;
  ram[2425]  = 93;
  ram[2426]  = 93;
  ram[2427]  = 94;
  ram[2428]  = 93;
  ram[2429]  = 93;
  ram[2430]  = 91;
  ram[2431]  = 92;
  ram[2432]  = 91;
  ram[2433]  = 92;
  ram[2434]  = 93;
  ram[2435]  = 93;
  ram[2436]  = 94;
  ram[2437]  = 93;
  ram[2438]  = 92;
  ram[2439]  = 91;
  ram[2440]  = 91;
  ram[2441]  = 91;
  ram[2442]  = 91;
  ram[2443]  = 92;
  ram[2444]  = 92;
  ram[2445]  = 91;
  ram[2446]  = 91;
  ram[2447]  = 92;
  ram[2448]  = 90;
  ram[2449]  = 90;
  ram[2450]  = 90;
  ram[2451]  = 90;
  ram[2452]  = 90;
  ram[2453]  = 91;
  ram[2454]  = 91;
  ram[2455]  = 91;
  ram[2456]  = 89;
  ram[2457]  = 90;
  ram[2458]  = 89;
  ram[2459]  = 90;
  ram[2460]  = 90;
  ram[2461]  = 91;
  ram[2462]  = 91;
  ram[2463]  = 91;
  ram[2464]  = 90;
  ram[2465]  = 89;
  ram[2466]  = 89;
  ram[2467]  = 91;
  ram[2468]  = 92;
  ram[2469]  = 91;
  ram[2470]  = 91;
  ram[2471]  = 90;
  ram[2472]  = 88;
  ram[2473]  = 89;
  ram[2474]  = 89;
  ram[2475]  = 91;
  ram[2476]  = 91;
  ram[2477]  = 91;
  ram[2478]  = 90;
  ram[2479]  = 90;
  ram[2480]  = 88;
  ram[2481]  = 90;
  ram[2482]  = 92;
  ram[2483]  = 92;
  ram[2484]  = 92;
  ram[2485]  = 91;
  ram[2486]  = 92;
  ram[2487]  = 92;
  ram[2488]  = 91;
  ram[2489]  = 91;
  ram[2490]  = 91;
  ram[2491]  = 92;
  ram[2492]  = 91;
  ram[2493]  = 91;
  ram[2494]  = 89;
  ram[2495]  = 90;
  ram[2496]  = 90;
  ram[2497]  = 90;
  ram[2498]  = 91;
  ram[2499]  = 91;
  ram[2500]  = 91;
  ram[2501]  = 90;
  ram[2502]  = 88;
  ram[2503]  = 87;
  ram[2504]  = 89;
  ram[2505]  = 88;
  ram[2506]  = 88;
  ram[2507]  = 89;
  ram[2508]  = 89;
  ram[2509]  = 89;
  ram[2510]  = 88;
  ram[2511]  = 89;
  ram[2512]  = 87;
  ram[2513]  = 86;
  ram[2514]  = 86;
  ram[2515]  = 87;
  ram[2516]  = 87;
  ram[2517]  = 87;
  ram[2518]  = 87;
  ram[2519]  = 89;
  ram[2520]  = 88;
  ram[2521]  = 88;
  ram[2522]  = 88;
  ram[2523]  = 89;
  ram[2524]  = 89;
  ram[2525]  = 89;
  ram[2526]  = 90;
  ram[2527]  = 90;
  ram[2528]  = 88;
  ram[2529]  = 87;
  ram[2530]  = 89;
  ram[2531]  = 90;
  ram[2532]  = 91;
  ram[2533]  = 90;
  ram[2534]  = 90;
  ram[2535]  = 89;
  ram[2536]  = 89;
  ram[2537]  = 88;
  ram[2538]  = 88;
  ram[2539]  = 89;
  ram[2540]  = 90;
  ram[2541]  = 89;
  ram[2542]  = 86;
  ram[2543]  = 86;
  ram[2544]  = 84;
  ram[2545]  = 86;
  ram[2546]  = 87;
  ram[2547]  = 88;
  ram[2548]  = 89;
  ram[2549]  = 89;
  ram[2550]  = 89;
  ram[2551]  = 90;
  ram[2552]  = 87;
  ram[2553]  = 88;
  ram[2554]  = 88;
  ram[2555]  = 88;
  ram[2556]  = 88;
  ram[2557]  = 87;
  ram[2558]  = 86;
  ram[2559]  = 86;
  ram[2560]  = 88;
  ram[2561]  = 88;
  ram[2562]  = 88;
  ram[2563]  = 87;
  ram[2564]  = 87;
  ram[2565]  = 87;
  ram[2566]  = 86;
  ram[2567]  = 86;
  ram[2568]  = 85;
  ram[2569]  = 86;
  ram[2570]  = 86;
  ram[2571]  = 85;
  ram[2572]  = 85;
  ram[2573]  = 85;
  ram[2574]  = 85;
  ram[2575]  = 87;
  ram[2576]  = 87;
  ram[2577]  = 73;
  ram[2578]  = 74;
  ram[2579]  = 72;
  ram[2580]  = 71;
  ram[2581]  = 72;
  ram[2582]  = 76;
  ram[2583]  = 73;
  ram[2584]  = 72;
  ram[2585]  = 74;
  ram[2586]  = 75;
  ram[2587]  = 72;
  ram[2588]  = 75;
  ram[2589]  = 74;
  ram[2590]  = 75;
  ram[2591]  = 76;
  ram[2592]  = 73;
  ram[2593]  = 71;
  ram[2594]  = 77;
  ram[2595]  = 73;
  ram[2596]  = 78;
  ram[2597]  = 77;
  ram[2598]  = 71;
  ram[2599]  = 78;
  ram[2600]  = 73;
  ram[2601]  = 74;
  ram[2602]  = 76;
  ram[2603]  = 73;
  ram[2604]  = 78;
  ram[2605]  = 80;
  ram[2606]  = 67;
  ram[2607]  = 85;
  ram[2608]  = 85;
  ram[2609]  = 86;
  ram[2610]  = 86;
  ram[2611]  = 85;
  ram[2612]  = 85;
  ram[2613]  = 85;
  ram[2614]  = 86;
  ram[2615]  = 86;
  ram[2616]  = 85;
  ram[2617]  = 87;
  ram[2618]  = 86;
  ram[2619]  = 86;
  ram[2620]  = 86;
  ram[2621]  = 85;
  ram[2622]  = 84;
  ram[2623]  = 83;
  ram[2624]  = 86;
  ram[2625]  = 86;
  ram[2626]  = 86;
  ram[2627]  = 86;
  ram[2628]  = 85;
  ram[2629]  = 85;
  ram[2630]  = 85;
  ram[2631]  = 85;
  ram[2632]  = 85;
  ram[2633]  = 85;
  ram[2634]  = 84;
  ram[2635]  = 84;
  ram[2636]  = 84;
  ram[2637]  = 84;
  ram[2638]  = 84;
  ram[2639]  = 85;
  ram[2640]  = 88;
  ram[2641]  = 177;
  ram[2642]  = 172;
  ram[2643]  = 175;
  ram[2644]  = 176;
  ram[2645]  = 172;
  ram[2646]  = 168;
  ram[2647]  = 176;
  ram[2648]  = 173;
  ram[2649]  = 176;
  ram[2650]  = 169;
  ram[2651]  = 176;
  ram[2652]  = 170;
  ram[2653]  = 178;
  ram[2654]  = 171;
  ram[2655]  = 174;
  ram[2656]  = 174;
  ram[2657]  = 177;
  ram[2658]  = 177;
  ram[2659]  = 172;
  ram[2660]  = 178;
  ram[2661]  = 168;
  ram[2662]  = 184;
  ram[2663]  = 169;
  ram[2664]  = 178;
  ram[2665]  = 175;
  ram[2666]  = 172;
  ram[2667]  = 173;
  ram[2668]  = 177;
  ram[2669]  = 168;
  ram[2670]  = 182;
  ram[2671]  = 89;
  ram[2672]  = 86;
  ram[2673]  = 87;
  ram[2674]  = 86;
  ram[2675]  = 84;
  ram[2676]  = 83;
  ram[2677]  = 84;
  ram[2678]  = 83;
  ram[2679]  = 83;
  ram[2680]  = 84;
  ram[2681]  = 84;
  ram[2682]  = 84;
  ram[2683]  = 84;
  ram[2684]  = 84;
  ram[2685]  = 84;
  ram[2686]  = 83;
  ram[2687]  = 83;
  ram[2688]  = 83;
  ram[2689]  = 83;
  ram[2690]  = 83;
  ram[2691]  = 82;
  ram[2692]  = 82;
  ram[2693]  = 82;
  ram[2694]  = 82;
  ram[2695]  = 82;
  ram[2696]  = 82;
  ram[2697]  = 81;
  ram[2698]  = 80;
  ram[2699]  = 81;
  ram[2700]  = 81;
  ram[2701]  = 81;
  ram[2702]  = 81;
  ram[2703]  = 82;
  ram[2704]  = 92;
  ram[2705]  = 248;
  ram[2706]  = 253;
  ram[2707]  = 247;
  ram[2708]  = 244;
  ram[2709]  = 250;
  ram[2710]  = 250;
  ram[2711]  = 249;
  ram[2712]  = 248;
  ram[2713]  = 249;
  ram[2714]  = 245;
  ram[2715]  = 250;
  ram[2716]  = 247;
  ram[2717]  = 251;
  ram[2718]  = 247;
  ram[2719]  = 247;
  ram[2720]  = 249;
  ram[2721]  = 245;
  ram[2722]  = 250;
  ram[2723]  = 248;
  ram[2724]  = 248;
  ram[2725]  = 248;
  ram[2726]  = 249;
  ram[2727]  = 253;
  ram[2728]  = 250;
  ram[2729]  = 246;
  ram[2730]  = 249;
  ram[2731]  = 251;
  ram[2732]  = 247;
  ram[2733]  = 237;
  ram[2734]  = 230;
  ram[2735]  = 95;
  ram[2736]  = 83;
  ram[2737]  = 82;
  ram[2738]  = 82;
  ram[2739]  = 82;
  ram[2740]  = 81;
  ram[2741]  = 81;
  ram[2742]  = 81;
  ram[2743]  = 82;
  ram[2744]  = 82;
  ram[2745]  = 81;
  ram[2746]  = 80;
  ram[2747]  = 81;
  ram[2748]  = 80;
  ram[2749]  = 81;
  ram[2750]  = 81;
  ram[2751]  = 82;
  ram[2752]  = 79;
  ram[2753]  = 79;
  ram[2754]  = 79;
  ram[2755]  = 79;
  ram[2756]  = 79;
  ram[2757]  = 78;
  ram[2758]  = 78;
  ram[2759]  = 78;
  ram[2760]  = 78;
  ram[2761]  = 78;
  ram[2762]  = 77;
  ram[2763]  = 78;
  ram[2764]  = 78;
  ram[2765]  = 79;
  ram[2766]  = 78;
  ram[2767]  = 79;
  ram[2768]  = 78;
  ram[2769]  = 114;
  ram[2770]  = 102;
  ram[2771]  = 106;
  ram[2772]  = 111;
  ram[2773]  = 104;
  ram[2774]  = 107;
  ram[2775]  = 108;
  ram[2776]  = 104;
  ram[2777]  = 108;
  ram[2778]  = 99;
  ram[2779]  = 114;
  ram[2780]  = 100;
  ram[2781]  = 112;
  ram[2782]  = 101;
  ram[2783]  = 103;
  ram[2784]  = 102;
  ram[2785]  = 110;
  ram[2786]  = 104;
  ram[2787]  = 100;
  ram[2788]  = 111;
  ram[2789]  = 101;
  ram[2790]  = 108;
  ram[2791]  = 102;
  ram[2792]  = 112;
  ram[2793]  = 103;
  ram[2794]  = 111;
  ram[2795]  = 99;
  ram[2796]  = 106;
  ram[2797]  = 212;
  ram[2798]  = 226;
  ram[2799]  = 87;
  ram[2800]  = 77;
  ram[2801]  = 77;
  ram[2802]  = 79;
  ram[2803]  = 78;
  ram[2804]  = 77;
  ram[2805]  = 78;
  ram[2806]  = 79;
  ram[2807]  = 80;
  ram[2808]  = 79;
  ram[2809]  = 79;
  ram[2810]  = 77;
  ram[2811]  = 78;
  ram[2812]  = 77;
  ram[2813]  = 78;
  ram[2814]  = 77;
  ram[2815]  = 79;
  ram[2816]  = 78;
  ram[2817]  = 78;
  ram[2818]  = 78;
  ram[2819]  = 77;
  ram[2820]  = 77;
  ram[2821]  = 77;
  ram[2822]  = 77;
  ram[2823]  = 77;
  ram[2824]  = 76;
  ram[2825]  = 77;
  ram[2826]  = 76;
  ram[2827]  = 77;
  ram[2828]  = 76;
  ram[2829]  = 76;
  ram[2830]  = 75;
  ram[2831]  = 76;
  ram[2832]  = 76;
  ram[2833]  = 62;
  ram[2834]  = 69;
  ram[2835]  = 66;
  ram[2836]  = 64;
  ram[2837]  = 60;
  ram[2838]  = 67;
  ram[2839]  = 64;
  ram[2840]  = 65;
  ram[2841]  = 63;
  ram[2842]  = 67;
  ram[2843]  = 65;
  ram[2844]  = 65;
  ram[2845]  = 62;
  ram[2846]  = 66;
  ram[2847]  = 62;
  ram[2848]  = 68;
  ram[2849]  = 61;
  ram[2850]  = 65;
  ram[2851]  = 67;
  ram[2852]  = 65;
  ram[2853]  = 66;
  ram[2854]  = 68;
  ram[2855]  = 61;
  ram[2856]  = 65;
  ram[2857]  = 67;
  ram[2858]  = 62;
  ram[2859]  = 62;
  ram[2860]  = 56;
  ram[2861]  = 215;
  ram[2862]  = 221;
  ram[2863]  = 84;
  ram[2864]  = 75;
  ram[2865]  = 76;
  ram[2866]  = 78;
  ram[2867]  = 77;
  ram[2868]  = 76;
  ram[2869]  = 76;
  ram[2870]  = 77;
  ram[2871]  = 77;
  ram[2872]  = 76;
  ram[2873]  = 76;
  ram[2874]  = 76;
  ram[2875]  = 77;
  ram[2876]  = 76;
  ram[2877]  = 76;
  ram[2878]  = 74;
  ram[2879]  = 75;
  ram[2880]  = 77;
  ram[2881]  = 78;
  ram[2882]  = 76;
  ram[2883]  = 77;
  ram[2884]  = 76;
  ram[2885]  = 76;
  ram[2886]  = 76;
  ram[2887]  = 76;
  ram[2888]  = 77;
  ram[2889]  = 78;
  ram[2890]  = 77;
  ram[2891]  = 77;
  ram[2892]  = 75;
  ram[2893]  = 75;
  ram[2894]  = 74;
  ram[2895]  = 74;
  ram[2896]  = 75;
  ram[2897]  = 70;
  ram[2898]  = 74;
  ram[2899]  = 70;
  ram[2900]  = 74;
  ram[2901]  = 72;
  ram[2902]  = 72;
  ram[2903]  = 71;
  ram[2904]  = 71;
  ram[2905]  = 71;
  ram[2906]  = 72;
  ram[2907]  = 75;
  ram[2908]  = 69;
  ram[2909]  = 76;
  ram[2910]  = 77;
  ram[2911]  = 72;
  ram[2912]  = 64;
  ram[2913]  = 67;
  ram[2914]  = 70;
  ram[2915]  = 74;
  ram[2916]  = 73;
  ram[2917]  = 70;
  ram[2918]  = 70;
  ram[2919]  = 71;
  ram[2920]  = 73;
  ram[2921]  = 70;
  ram[2922]  = 71;
  ram[2923]  = 61;
  ram[2924]  = 65;
  ram[2925]  = 209;
  ram[2926]  = 218;
  ram[2927]  = 81;
  ram[2928]  = 75;
  ram[2929]  = 75;
  ram[2930]  = 77;
  ram[2931]  = 76;
  ram[2932]  = 76;
  ram[2933]  = 76;
  ram[2934]  = 77;
  ram[2935]  = 77;
  ram[2936]  = 76;
  ram[2937]  = 76;
  ram[2938]  = 76;
  ram[2939]  = 77;
  ram[2940]  = 76;
  ram[2941]  = 76;
  ram[2942]  = 74;
  ram[2943]  = 75;
  ram[2944]  = 75;
  ram[2945]  = 76;
  ram[2946]  = 75;
  ram[2947]  = 75;
  ram[2948]  = 75;
  ram[2949]  = 75;
  ram[2950]  = 74;
  ram[2951]  = 74;
  ram[2952]  = 76;
  ram[2953]  = 75;
  ram[2954]  = 74;
  ram[2955]  = 74;
  ram[2956]  = 73;
  ram[2957]  = 73;
  ram[2958]  = 72;
  ram[2959]  = 72;
  ram[2960]  = 72;
  ram[2961]  = 80;
  ram[2962]  = 76;
  ram[2963]  = 74;
  ram[2964]  = 76;
  ram[2965]  = 74;
  ram[2966]  = 70;
  ram[2967]  = 70;
  ram[2968]  = 73;
  ram[2969]  = 69;
  ram[2970]  = 74;
  ram[2971]  = 69;
  ram[2972]  = 74;
  ram[2973]  = 75;
  ram[2974]  = 77;
  ram[2975]  = 63;
  ram[2976]  = 85;
  ram[2977]  = 79;
  ram[2978]  = 66;
  ram[2979]  = 74;
  ram[2980]  = 72;
  ram[2981]  = 75;
  ram[2982]  = 71;
  ram[2983]  = 76;
  ram[2984]  = 87;
  ram[2985]  = 82;
  ram[2986]  = 79;
  ram[2987]  = 84;
  ram[2988]  = 73;
  ram[2989]  = 218;
  ram[2990]  = 228;
  ram[2991]  = 75;
  ram[2992]  = 73;
  ram[2993]  = 72;
  ram[2994]  = 74;
  ram[2995]  = 74;
  ram[2996]  = 75;
  ram[2997]  = 75;
  ram[2998]  = 76;
  ram[2999]  = 75;
  ram[3000]  = 75;
  ram[3001]  = 75;
  ram[3002]  = 74;
  ram[3003]  = 75;
  ram[3004]  = 74;
  ram[3005]  = 75;
  ram[3006]  = 73;
  ram[3007]  = 74;
  ram[3008]  = 73;
  ram[3009]  = 73;
  ram[3010]  = 72;
  ram[3011]  = 73;
  ram[3012]  = 72;
  ram[3013]  = 72;
  ram[3014]  = 72;
  ram[3015]  = 72;
  ram[3016]  = 72;
  ram[3017]  = 71;
  ram[3018]  = 71;
  ram[3019]  = 70;
  ram[3020]  = 70;
  ram[3021]  = 71;
  ram[3022]  = 71;
  ram[3023]  = 71;
  ram[3024]  = 74;
  ram[3025]  = 73;
  ram[3026]  = 71;
  ram[3027]  = 75;
  ram[3028]  = 72;
  ram[3029]  = 72;
  ram[3030]  = 71;
  ram[3031]  = 72;
  ram[3032]  = 73;
  ram[3033]  = 70;
  ram[3034]  = 71;
  ram[3035]  = 71;
  ram[3036]  = 71;
  ram[3037]  = 74;
  ram[3038]  = 66;
  ram[3039]  = 46;
  ram[3040]  = 255;
  ram[3041]  = 255;
  ram[3042]  = 41;
  ram[3043]  = 72;
  ram[3044]  = 75;
  ram[3045]  = 71;
  ram[3046]  = 61;
  ram[3047]  = 163;
  ram[3048]  = 241;
  ram[3049]  = 219;
  ram[3050]  = 225;
  ram[3051]  = 224;
  ram[3052]  = 226;
  ram[3053]  = 216;
  ram[3054]  = 225;
  ram[3055]  = 82;
  ram[3056]  = 73;
  ram[3057]  = 71;
  ram[3058]  = 72;
  ram[3059]  = 72;
  ram[3060]  = 72;
  ram[3061]  = 72;
  ram[3062]  = 71;
  ram[3063]  = 70;
  ram[3064]  = 71;
  ram[3065]  = 71;
  ram[3066]  = 71;
  ram[3067]  = 71;
  ram[3068]  = 71;
  ram[3069]  = 71;
  ram[3070]  = 72;
  ram[3071]  = 72;
  ram[3072]  = 69;
  ram[3073]  = 70;
  ram[3074]  = 70;
  ram[3075]  = 71;
  ram[3076]  = 71;
  ram[3077]  = 71;
  ram[3078]  = 70;
  ram[3079]  = 70;
  ram[3080]  = 71;
  ram[3081]  = 71;
  ram[3082]  = 71;
  ram[3083]  = 70;
  ram[3084]  = 70;
  ram[3085]  = 70;
  ram[3086]  = 70;
  ram[3087]  = 71;
  ram[3088]  = 69;
  ram[3089]  = 68;
  ram[3090]  = 67;
  ram[3091]  = 68;
  ram[3092]  = 69;
  ram[3093]  = 70;
  ram[3094]  = 69;
  ram[3095]  = 67;
  ram[3096]  = 70;
  ram[3097]  = 69;
  ram[3098]  = 69;
  ram[3099]  = 70;
  ram[3100]  = 67;
  ram[3101]  = 72;
  ram[3102]  = 69;
  ram[3103]  = 44;
  ram[3104]  = 239;
  ram[3105]  = 223;
  ram[3106]  = 39;
  ram[3107]  = 67;
  ram[3108]  = 70;
  ram[3109]  = 72;
  ram[3110]  = 59;
  ram[3111]  = 138;
  ram[3112]  = 214;
  ram[3113]  = 207;
  ram[3114]  = 205;
  ram[3115]  = 201;
  ram[3116]  = 205;
  ram[3117]  = 203;
  ram[3118]  = 193;
  ram[3119]  = 76;
  ram[3120]  = 71;
  ram[3121]  = 68;
  ram[3122]  = 68;
  ram[3123]  = 70;
  ram[3124]  = 69;
  ram[3125]  = 71;
  ram[3126]  = 71;
  ram[3127]  = 71;
  ram[3128]  = 71;
  ram[3129]  = 71;
  ram[3130]  = 71;
  ram[3131]  = 70;
  ram[3132]  = 70;
  ram[3133]  = 70;
  ram[3134]  = 69;
  ram[3135]  = 68;
  ram[3136]  = 70;
  ram[3137]  = 70;
  ram[3138]  = 70;
  ram[3139]  = 71;
  ram[3140]  = 71;
  ram[3141]  = 70;
  ram[3142]  = 70;
  ram[3143]  = 70;
  ram[3144]  = 69;
  ram[3145]  = 69;
  ram[3146]  = 69;
  ram[3147]  = 69;
  ram[3148]  = 69;
  ram[3149]  = 69;
  ram[3150]  = 70;
  ram[3151]  = 70;
  ram[3152]  = 68;
  ram[3153]  = 67;
  ram[3154]  = 67;
  ram[3155]  = 67;
  ram[3156]  = 69;
  ram[3157]  = 69;
  ram[3158]  = 68;
  ram[3159]  = 67;
  ram[3160]  = 67;
  ram[3161]  = 67;
  ram[3162]  = 68;
  ram[3163]  = 70;
  ram[3164]  = 66;
  ram[3165]  = 68;
  ram[3166]  = 71;
  ram[3167]  = 59;
  ram[3168]  = 65;
  ram[3169]  = 58;
  ram[3170]  = 67;
  ram[3171]  = 69;
  ram[3172]  = 68;
  ram[3173]  = 74;
  ram[3174]  = 69;
  ram[3175]  = 68;
  ram[3176]  = 58;
  ram[3177]  = 61;
  ram[3178]  = 64;
  ram[3179]  = 59;
  ram[3180]  = 66;
  ram[3181]  = 57;
  ram[3182]  = 65;
  ram[3183]  = 67;
  ram[3184]  = 69;
  ram[3185]  = 68;
  ram[3186]  = 70;
  ram[3187]  = 70;
  ram[3188]  = 70;
  ram[3189]  = 71;
  ram[3190]  = 70;
  ram[3191]  = 70;
  ram[3192]  = 69;
  ram[3193]  = 70;
  ram[3194]  = 70;
  ram[3195]  = 69;
  ram[3196]  = 69;
  ram[3197]  = 69;
  ram[3198]  = 68;
  ram[3199]  = 67;
  ram[3200]  = 69;
  ram[3201]  = 69;
  ram[3202]  = 69;
  ram[3203]  = 69;
  ram[3204]  = 69;
  ram[3205]  = 68;
  ram[3206]  = 68;
  ram[3207]  = 68;
  ram[3208]  = 68;
  ram[3209]  = 67;
  ram[3210]  = 67;
  ram[3211]  = 67;
  ram[3212]  = 68;
  ram[3213]  = 68;
  ram[3214]  = 68;
  ram[3215]  = 68;
  ram[3216]  = 68;
  ram[3217]  = 67;
  ram[3218]  = 67;
  ram[3219]  = 67;
  ram[3220]  = 68;
  ram[3221]  = 69;
  ram[3222]  = 68;
  ram[3223]  = 67;
  ram[3224]  = 66;
  ram[3225]  = 66;
  ram[3226]  = 67;
  ram[3227]  = 69;
  ram[3228]  = 67;
  ram[3229]  = 66;
  ram[3230]  = 71;
  ram[3231]  = 69;
  ram[3232]  = 59;
  ram[3233]  = 66;
  ram[3234]  = 66;
  ram[3235]  = 70;
  ram[3236]  = 73;
  ram[3237]  = 68;
  ram[3238]  = 69;
  ram[3239]  = 66;
  ram[3240]  = 72;
  ram[3241]  = 66;
  ram[3242]  = 68;
  ram[3243]  = 63;
  ram[3244]  = 61;
  ram[3245]  = 69;
  ram[3246]  = 66;
  ram[3247]  = 71;
  ram[3248]  = 68;
  ram[3249]  = 68;
  ram[3250]  = 68;
  ram[3251]  = 68;
  ram[3252]  = 69;
  ram[3253]  = 69;
  ram[3254]  = 70;
  ram[3255]  = 70;
  ram[3256]  = 68;
  ram[3257]  = 69;
  ram[3258]  = 69;
  ram[3259]  = 68;
  ram[3260]  = 68;
  ram[3261]  = 68;
  ram[3262]  = 68;
  ram[3263]  = 67;
  ram[3264]  = 69;
  ram[3265]  = 69;
  ram[3266]  = 69;
  ram[3267]  = 69;
  ram[3268]  = 68;
  ram[3269]  = 68;
  ram[3270]  = 68;
  ram[3271]  = 68;
  ram[3272]  = 68;
  ram[3273]  = 68;
  ram[3274]  = 68;
  ram[3275]  = 68;
  ram[3276]  = 69;
  ram[3277]  = 69;
  ram[3278]  = 69;
  ram[3279]  = 69;
  ram[3280]  = 69;
  ram[3281]  = 68;
  ram[3282]  = 68;
  ram[3283]  = 68;
  ram[3284]  = 69;
  ram[3285]  = 69;
  ram[3286]  = 68;
  ram[3287]  = 67;
  ram[3288]  = 68;
  ram[3289]  = 68;
  ram[3290]  = 66;
  ram[3291]  = 68;
  ram[3292]  = 69;
  ram[3293]  = 68;
  ram[3294]  = 68;
  ram[3295]  = 68;
  ram[3296]  = 70;
  ram[3297]  = 68;
  ram[3298]  = 66;
  ram[3299]  = 74;
  ram[3300]  = 68;
  ram[3301]  = 70;
  ram[3302]  = 74;
  ram[3303]  = 71;
  ram[3304]  = 64;
  ram[3305]  = 69;
  ram[3306]  = 68;
  ram[3307]  = 70;
  ram[3308]  = 66;
  ram[3309]  = 68;
  ram[3310]  = 68;
  ram[3311]  = 70;
  ram[3312]  = 67;
  ram[3313]  = 68;
  ram[3314]  = 67;
  ram[3315]  = 69;
  ram[3316]  = 68;
  ram[3317]  = 70;
  ram[3318]  = 69;
  ram[3319]  = 70;
  ram[3320]  = 69;
  ram[3321]  = 70;
  ram[3322]  = 69;
  ram[3323]  = 69;
  ram[3324]  = 68;
  ram[3325]  = 68;
  ram[3326]  = 68;
  ram[3327]  = 67;
  ram[3328]  = 70;
  ram[3329]  = 70;
  ram[3330]  = 70;
  ram[3331]  = 70;
  ram[3332]  = 70;
  ram[3333]  = 70;
  ram[3334]  = 70;
  ram[3335]  = 70;
  ram[3336]  = 70;
  ram[3337]  = 70;
  ram[3338]  = 70;
  ram[3339]  = 70;
  ram[3340]  = 70;
  ram[3341]  = 70;
  ram[3342]  = 70;
  ram[3343]  = 70;
  ram[3344]  = 69;
  ram[3345]  = 69;
  ram[3346]  = 68;
  ram[3347]  = 69;
  ram[3348]  = 69;
  ram[3349]  = 69;
  ram[3350]  = 69;
  ram[3351]  = 68;
  ram[3352]  = 68;
  ram[3353]  = 70;
  ram[3354]  = 68;
  ram[3355]  = 67;
  ram[3356]  = 69;
  ram[3357]  = 69;
  ram[3358]  = 67;
  ram[3359]  = 67;
  ram[3360]  = 67;
  ram[3361]  = 68;
  ram[3362]  = 72;
  ram[3363]  = 68;
  ram[3364]  = 69;
  ram[3365]  = 75;
  ram[3366]  = 68;
  ram[3367]  = 72;
  ram[3368]  = 72;
  ram[3369]  = 67;
  ram[3370]  = 65;
  ram[3371]  = 72;
  ram[3372]  = 70;
  ram[3373]  = 65;
  ram[3374]  = 72;
  ram[3375]  = 69;
  ram[3376]  = 69;
  ram[3377]  = 69;
  ram[3378]  = 68;
  ram[3379]  = 70;
  ram[3380]  = 69;
  ram[3381]  = 70;
  ram[3382]  = 69;
  ram[3383]  = 71;
  ram[3384]  = 70;
  ram[3385]  = 70;
  ram[3386]  = 70;
  ram[3387]  = 69;
  ram[3388]  = 69;
  ram[3389]  = 69;
  ram[3390]  = 68;
  ram[3391]  = 67;
  ram[3392]  = 70;
  ram[3393]  = 70;
  ram[3394]  = 70;
  ram[3395]  = 70;
  ram[3396]  = 70;
  ram[3397]  = 71;
  ram[3398]  = 71;
  ram[3399]  = 71;
  ram[3400]  = 72;
  ram[3401]  = 72;
  ram[3402]  = 72;
  ram[3403]  = 72;
  ram[3404]  = 72;
  ram[3405]  = 72;
  ram[3406]  = 72;
  ram[3407]  = 71;
  ram[3408]  = 69;
  ram[3409]  = 69;
  ram[3410]  = 68;
  ram[3411]  = 69;
  ram[3412]  = 69;
  ram[3413]  = 69;
  ram[3414]  = 68;
  ram[3415]  = 68;
  ram[3416]  = 66;
  ram[3417]  = 69;
  ram[3418]  = 71;
  ram[3419]  = 67;
  ram[3420]  = 67;
  ram[3421]  = 69;
  ram[3422]  = 68;
  ram[3423]  = 71;
  ram[3424]  = 73;
  ram[3425]  = 68;
  ram[3426]  = 65;
  ram[3427]  = 77;
  ram[3428]  = 69;
  ram[3429]  = 72;
  ram[3430]  = 74;
  ram[3431]  = 70;
  ram[3432]  = 66;
  ram[3433]  = 74;
  ram[3434]  = 73;
  ram[3435]  = 65;
  ram[3436]  = 74;
  ram[3437]  = 68;
  ram[3438]  = 66;
  ram[3439]  = 75;
  ram[3440]  = 72;
  ram[3441]  = 70;
  ram[3442]  = 70;
  ram[3443]  = 69;
  ram[3444]  = 69;
  ram[3445]  = 69;
  ram[3446]  = 69;
  ram[3447]  = 69;
  ram[3448]  = 71;
  ram[3449]  = 72;
  ram[3450]  = 72;
  ram[3451]  = 71;
  ram[3452]  = 70;
  ram[3453]  = 70;
  ram[3454]  = 69;
  ram[3455]  = 68;
  ram[3456]  = 69;
  ram[3457]  = 69;
  ram[3458]  = 69;
  ram[3459]  = 69;
  ram[3460]  = 70;
  ram[3461]  = 70;
  ram[3462]  = 71;
  ram[3463]  = 71;
  ram[3464]  = 72;
  ram[3465]  = 72;
  ram[3466]  = 72;
  ram[3467]  = 72;
  ram[3468]  = 72;
  ram[3469]  = 71;
  ram[3470]  = 71;
  ram[3471]  = 70;
  ram[3472]  = 69;
  ram[3473]  = 69;
  ram[3474]  = 68;
  ram[3475]  = 68;
  ram[3476]  = 69;
  ram[3477]  = 68;
  ram[3478]  = 68;
  ram[3479]  = 67;
  ram[3480]  = 67;
  ram[3481]  = 67;
  ram[3482]  = 71;
  ram[3483]  = 69;
  ram[3484]  = 67;
  ram[3485]  = 70;
  ram[3486]  = 69;
  ram[3487]  = 72;
  ram[3488]  = 67;
  ram[3489]  = 66;
  ram[3490]  = 75;
  ram[3491]  = 71;
  ram[3492]  = 66;
  ram[3493]  = 69;
  ram[3494]  = 74;
  ram[3495]  = 69;
  ram[3496]  = 80;
  ram[3497]  = 67;
  ram[3498]  = 71;
  ram[3499]  = 71;
  ram[3500]  = 68;
  ram[3501]  = 68;
  ram[3502]  = 71;
  ram[3503]  = 70;
  ram[3504]  = 71;
  ram[3505]  = 69;
  ram[3506]  = 69;
  ram[3507]  = 69;
  ram[3508]  = 69;
  ram[3509]  = 69;
  ram[3510]  = 69;
  ram[3511]  = 69;
  ram[3512]  = 71;
  ram[3513]  = 72;
  ram[3514]  = 72;
  ram[3515]  = 71;
  ram[3516]  = 70;
  ram[3517]  = 70;
  ram[3518]  = 69;
  ram[3519]  = 68;
  ram[3520]  = 71;
  ram[3521]  = 70;
  ram[3522]  = 70;
  ram[3523]  = 71;
  ram[3524]  = 71;
  ram[3525]  = 72;
  ram[3526]  = 72;
  ram[3527]  = 73;
  ram[3528]  = 72;
  ram[3529]  = 72;
  ram[3530]  = 72;
  ram[3531]  = 72;
  ram[3532]  = 72;
  ram[3533]  = 71;
  ram[3534]  = 70;
  ram[3535]  = 70;
  ram[3536]  = 71;
  ram[3537]  = 70;
  ram[3538]  = 70;
  ram[3539]  = 70;
  ram[3540]  = 70;
  ram[3541]  = 70;
  ram[3542]  = 69;
  ram[3543]  = 69;
  ram[3544]  = 71;
  ram[3545]  = 67;
  ram[3546]  = 72;
  ram[3547]  = 72;
  ram[3548]  = 72;
  ram[3549]  = 73;
  ram[3550]  = 70;
  ram[3551]  = 70;
  ram[3552]  = 70;
  ram[3553]  = 75;
  ram[3554]  = 66;
  ram[3555]  = 72;
  ram[3556]  = 72;
  ram[3557]  = 70;
  ram[3558]  = 68;
  ram[3559]  = 70;
  ram[3560]  = 70;
  ram[3561]  = 76;
  ram[3562]  = 71;
  ram[3563]  = 69;
  ram[3564]  = 70;
  ram[3565]  = 73;
  ram[3566]  = 71;
  ram[3567]  = 67;
  ram[3568]  = 70;
  ram[3569]  = 70;
  ram[3570]  = 70;
  ram[3571]  = 70;
  ram[3572]  = 71;
  ram[3573]  = 71;
  ram[3574]  = 71;
  ram[3575]  = 72;
  ram[3576]  = 71;
  ram[3577]  = 72;
  ram[3578]  = 73;
  ram[3579]  = 72;
  ram[3580]  = 71;
  ram[3581]  = 71;
  ram[3582]  = 70;
  ram[3583]  = 68;
  ram[3584]  = 72;
  ram[3585]  = 72;
  ram[3586]  = 72;
  ram[3587]  = 71;
  ram[3588]  = 71;
  ram[3589]  = 71;
  ram[3590]  = 71;
  ram[3591]  = 70;
  ram[3592]  = 70;
  ram[3593]  = 70;
  ram[3594]  = 70;
  ram[3595]  = 70;
  ram[3596]  = 70;
  ram[3597]  = 70;
  ram[3598]  = 70;
  ram[3599]  = 70;
  ram[3600]  = 69;
  ram[3601]  = 69;
  ram[3602]  = 69;
  ram[3603]  = 70;
  ram[3604]  = 70;
  ram[3605]  = 70;
  ram[3606]  = 70;
  ram[3607]  = 70;
  ram[3608]  = 70;
  ram[3609]  = 70;
  ram[3610]  = 70;
  ram[3611]  = 70;
  ram[3612]  = 70;
  ram[3613]  = 70;
  ram[3614]  = 70;
  ram[3615]  = 70;
  ram[3616]  = 71;
  ram[3617]  = 72;
  ram[3618]  = 71;
  ram[3619]  = 71;
  ram[3620]  = 71;
  ram[3621]  = 71;
  ram[3622]  = 71;
  ram[3623]  = 71;
  ram[3624]  = 70;
  ram[3625]  = 70;
  ram[3626]  = 70;
  ram[3627]  = 70;
  ram[3628]  = 70;
  ram[3629]  = 70;
  ram[3630]  = 70;
  ram[3631]  = 70;
  ram[3632]  = 71;
  ram[3633]  = 71;
  ram[3634]  = 71;
  ram[3635]  = 71;
  ram[3636]  = 71;
  ram[3637]  = 71;
  ram[3638]  = 71;
  ram[3639]  = 71;
  ram[3640]  = 72;
  ram[3641]  = 72;
  ram[3642]  = 72;
  ram[3643]  = 72;
  ram[3644]  = 71;
  ram[3645]  = 70;
  ram[3646]  = 70;
  ram[3647]  = 69;
  ram[3648]  = 71;
  ram[3649]  = 72;
  ram[3650]  = 72;
  ram[3651]  = 71;
  ram[3652]  = 71;
  ram[3653]  = 72;
  ram[3654]  = 72;
  ram[3655]  = 71;
  ram[3656]  = 73;
  ram[3657]  = 73;
  ram[3658]  = 73;
  ram[3659]  = 73;
  ram[3660]  = 73;
  ram[3661]  = 73;
  ram[3662]  = 73;
  ram[3663]  = 73;
  ram[3664]  = 73;
  ram[3665]  = 73;
  ram[3666]  = 73;
  ram[3667]  = 73;
  ram[3668]  = 73;
  ram[3669]  = 73;
  ram[3670]  = 73;
  ram[3671]  = 73;
  ram[3672]  = 72;
  ram[3673]  = 72;
  ram[3674]  = 72;
  ram[3675]  = 72;
  ram[3676]  = 72;
  ram[3677]  = 72;
  ram[3678]  = 72;
  ram[3679]  = 72;
  ram[3680]  = 73;
  ram[3681]  = 73;
  ram[3682]  = 73;
  ram[3683]  = 73;
  ram[3684]  = 73;
  ram[3685]  = 73;
  ram[3686]  = 72;
  ram[3687]  = 72;
  ram[3688]  = 72;
  ram[3689]  = 72;
  ram[3690]  = 71;
  ram[3691]  = 71;
  ram[3692]  = 71;
  ram[3693]  = 71;
  ram[3694]  = 72;
  ram[3695]  = 72;
  ram[3696]  = 72;
  ram[3697]  = 72;
  ram[3698]  = 72;
  ram[3699]  = 72;
  ram[3700]  = 73;
  ram[3701]  = 73;
  ram[3702]  = 73;
  ram[3703]  = 73;
  ram[3704]  = 72;
  ram[3705]  = 72;
  ram[3706]  = 72;
  ram[3707]  = 72;
  ram[3708]  = 71;
  ram[3709]  = 70;
  ram[3710]  = 70;
  ram[3711]  = 69;
  ram[3712]  = 72;
  ram[3713]  = 72;
  ram[3714]  = 72;
  ram[3715]  = 71;
  ram[3716]  = 72;
  ram[3717]  = 73;
  ram[3718]  = 73;
  ram[3719]  = 73;
  ram[3720]  = 73;
  ram[3721]  = 73;
  ram[3722]  = 73;
  ram[3723]  = 73;
  ram[3724]  = 72;
  ram[3725]  = 72;
  ram[3726]  = 72;
  ram[3727]  = 72;
  ram[3728]  = 72;
  ram[3729]  = 72;
  ram[3730]  = 72;
  ram[3731]  = 72;
  ram[3732]  = 72;
  ram[3733]  = 72;
  ram[3734]  = 72;
  ram[3735]  = 72;
  ram[3736]  = 72;
  ram[3737]  = 72;
  ram[3738]  = 72;
  ram[3739]  = 72;
  ram[3740]  = 72;
  ram[3741]  = 72;
  ram[3742]  = 72;
  ram[3743]  = 72;
  ram[3744]  = 73;
  ram[3745]  = 73;
  ram[3746]  = 73;
  ram[3747]  = 73;
  ram[3748]  = 73;
  ram[3749]  = 72;
  ram[3750]  = 72;
  ram[3751]  = 72;
  ram[3752]  = 73;
  ram[3753]  = 73;
  ram[3754]  = 73;
  ram[3755]  = 73;
  ram[3756]  = 72;
  ram[3757]  = 72;
  ram[3758]  = 72;
  ram[3759]  = 73;
  ram[3760]  = 71;
  ram[3761]  = 71;
  ram[3762]  = 71;
  ram[3763]  = 71;
  ram[3764]  = 72;
  ram[3765]  = 72;
  ram[3766]  = 72;
  ram[3767]  = 72;
  ram[3768]  = 72;
  ram[3769]  = 72;
  ram[3770]  = 72;
  ram[3771]  = 72;
  ram[3772]  = 71;
  ram[3773]  = 70;
  ram[3774]  = 70;
  ram[3775]  = 69;
  ram[3776]  = 73;
  ram[3777]  = 73;
  ram[3778]  = 73;
  ram[3779]  = 72;
  ram[3780]  = 72;
  ram[3781]  = 73;
  ram[3782]  = 73;
  ram[3783]  = 73;
  ram[3784]  = 74;
  ram[3785]  = 73;
  ram[3786]  = 73;
  ram[3787]  = 73;
  ram[3788]  = 73;
  ram[3789]  = 73;
  ram[3790]  = 73;
  ram[3791]  = 73;
  ram[3792]  = 73;
  ram[3793]  = 73;
  ram[3794]  = 73;
  ram[3795]  = 73;
  ram[3796]  = 73;
  ram[3797]  = 73;
  ram[3798]  = 73;
  ram[3799]  = 73;
  ram[3800]  = 74;
  ram[3801]  = 74;
  ram[3802]  = 74;
  ram[3803]  = 74;
  ram[3804]  = 74;
  ram[3805]  = 73;
  ram[3806]  = 73;
  ram[3807]  = 73;
  ram[3808]  = 75;
  ram[3809]  = 75;
  ram[3810]  = 75;
  ram[3811]  = 74;
  ram[3812]  = 74;
  ram[3813]  = 74;
  ram[3814]  = 74;
  ram[3815]  = 74;
  ram[3816]  = 75;
  ram[3817]  = 75;
  ram[3818]  = 74;
  ram[3819]  = 74;
  ram[3820]  = 74;
  ram[3821]  = 75;
  ram[3822]  = 74;
  ram[3823]  = 74;
  ram[3824]  = 74;
  ram[3825]  = 74;
  ram[3826]  = 72;
  ram[3827]  = 73;
  ram[3828]  = 73;
  ram[3829]  = 73;
  ram[3830]  = 73;
  ram[3831]  = 73;
  ram[3832]  = 72;
  ram[3833]  = 72;
  ram[3834]  = 72;
  ram[3835]  = 72;
  ram[3836]  = 71;
  ram[3837]  = 70;
  ram[3838]  = 70;
  ram[3839]  = 69;
  ram[3840]  = 74;
  ram[3841]  = 74;
  ram[3842]  = 73;
  ram[3843]  = 72;
  ram[3844]  = 72;
  ram[3845]  = 72;
  ram[3846]  = 72;
  ram[3847]  = 72;
  ram[3848]  = 72;
  ram[3849]  = 72;
  ram[3850]  = 72;
  ram[3851]  = 72;
  ram[3852]  = 72;
  ram[3853]  = 72;
  ram[3854]  = 72;
  ram[3855]  = 72;
  ram[3856]  = 73;
  ram[3857]  = 73;
  ram[3858]  = 73;
  ram[3859]  = 73;
  ram[3860]  = 73;
  ram[3861]  = 73;
  ram[3862]  = 74;
  ram[3863]  = 74;
  ram[3864]  = 73;
  ram[3865]  = 73;
  ram[3866]  = 73;
  ram[3867]  = 73;
  ram[3868]  = 73;
  ram[3869]  = 73;
  ram[3870]  = 73;
  ram[3871]  = 73;
  ram[3872]  = 73;
  ram[3873]  = 74;
  ram[3874]  = 73;
  ram[3875]  = 73;
  ram[3876]  = 73;
  ram[3877]  = 73;
  ram[3878]  = 73;
  ram[3879]  = 73;
  ram[3880]  = 73;
  ram[3881]  = 73;
  ram[3882]  = 73;
  ram[3883]  = 73;
  ram[3884]  = 73;
  ram[3885]  = 73;
  ram[3886]  = 72;
  ram[3887]  = 72;
  ram[3888]  = 73;
  ram[3889]  = 73;
  ram[3890]  = 72;
  ram[3891]  = 71;
  ram[3892]  = 71;
  ram[3893]  = 71;
  ram[3894]  = 71;
  ram[3895]  = 72;
  ram[3896]  = 72;
  ram[3897]  = 72;
  ram[3898]  = 72;
  ram[3899]  = 72;
  ram[3900]  = 71;
  ram[3901]  = 71;
  ram[3902]  = 70;
  ram[3903]  = 69;
  ram[3904]  = 73;
  ram[3905]  = 74;
  ram[3906]  = 73;
  ram[3907]  = 72;
  ram[3908]  = 71;
  ram[3909]  = 72;
  ram[3910]  = 72;
  ram[3911]  = 71;
  ram[3912]  = 71;
  ram[3913]  = 71;
  ram[3914]  = 71;
  ram[3915]  = 71;
  ram[3916]  = 71;
  ram[3917]  = 71;
  ram[3918]  = 71;
  ram[3919]  = 71;
  ram[3920]  = 71;
  ram[3921]  = 71;
  ram[3922]  = 71;
  ram[3923]  = 72;
  ram[3924]  = 72;
  ram[3925]  = 72;
  ram[3926]  = 72;
  ram[3927]  = 72;
  ram[3928]  = 72;
  ram[3929]  = 71;
  ram[3930]  = 71;
  ram[3931]  = 71;
  ram[3932]  = 71;
  ram[3933]  = 71;
  ram[3934]  = 71;
  ram[3935]  = 71;
  ram[3936]  = 72;
  ram[3937]  = 72;
  ram[3938]  = 71;
  ram[3939]  = 71;
  ram[3940]  = 71;
  ram[3941]  = 71;
  ram[3942]  = 71;
  ram[3943]  = 71;
  ram[3944]  = 71;
  ram[3945]  = 71;
  ram[3946]  = 71;
  ram[3947]  = 71;
  ram[3948]  = 71;
  ram[3949]  = 71;
  ram[3950]  = 70;
  ram[3951]  = 70;
  ram[3952]  = 71;
  ram[3953]  = 71;
  ram[3954]  = 71;
  ram[3955]  = 71;
  ram[3956]  = 70;
  ram[3957]  = 70;
  ram[3958]  = 70;
  ram[3959]  = 70;
  ram[3960]  = 72;
  ram[3961]  = 72;
  ram[3962]  = 72;
  ram[3963]  = 72;
  ram[3964]  = 71;
  ram[3965]  = 71;
  ram[3966]  = 70;
  ram[3967]  = 69;
  ram[3968]  = 71;
  ram[3969]  = 72;
  ram[3970]  = 72;
  ram[3971]  = 71;
  ram[3972]  = 71;
  ram[3973]  = 72;
  ram[3974]  = 72;
  ram[3975]  = 72;
  ram[3976]  = 74;
  ram[3977]  = 74;
  ram[3978]  = 74;
  ram[3979]  = 74;
  ram[3980]  = 74;
  ram[3981]  = 74;
  ram[3982]  = 74;
  ram[3983]  = 74;
  ram[3984]  = 73;
  ram[3985]  = 73;
  ram[3986]  = 74;
  ram[3987]  = 74;
  ram[3988]  = 74;
  ram[3989]  = 74;
  ram[3990]  = 74;
  ram[3991]  = 74;
  ram[3992]  = 74;
  ram[3993]  = 74;
  ram[3994]  = 74;
  ram[3995]  = 74;
  ram[3996]  = 74;
  ram[3997]  = 74;
  ram[3998]  = 74;
  ram[3999]  = 74;
  ram[4000]  = 74;
  ram[4001]  = 74;
  ram[4002]  = 74;
  ram[4003]  = 74;
  ram[4004]  = 73;
  ram[4005]  = 73;
  ram[4006]  = 73;
  ram[4007]  = 74;
  ram[4008]  = 74;
  ram[4009]  = 74;
  ram[4010]  = 74;
  ram[4011]  = 74;
  ram[4012]  = 73;
  ram[4013]  = 73;
  ram[4014]  = 74;
  ram[4015]  = 74;
  ram[4016]  = 74;
  ram[4017]  = 74;
  ram[4018]  = 74;
  ram[4019]  = 74;
  ram[4020]  = 74;
  ram[4021]  = 74;
  ram[4022]  = 74;
  ram[4023]  = 74;
  ram[4024]  = 73;
  ram[4025]  = 73;
  ram[4026]  = 72;
  ram[4027]  = 72;
  ram[4028]  = 71;
  ram[4029]  = 71;
  ram[4030]  = 70;
  ram[4031]  = 69;
  ram[4032]  = 69;
  ram[4033]  = 70;
  ram[4034]  = 71;
  ram[4035]  = 71;
  ram[4036]  = 72;
  ram[4037]  = 73;
  ram[4038]  = 73;
  ram[4039]  = 72;
  ram[4040]  = 71;
  ram[4041]  = 71;
  ram[4042]  = 71;
  ram[4043]  = 71;
  ram[4044]  = 71;
  ram[4045]  = 71;
  ram[4046]  = 71;
  ram[4047]  = 71;
  ram[4048]  = 72;
  ram[4049]  = 72;
  ram[4050]  = 72;
  ram[4051]  = 72;
  ram[4052]  = 72;
  ram[4053]  = 72;
  ram[4054]  = 72;
  ram[4055]  = 72;
  ram[4056]  = 72;
  ram[4057]  = 72;
  ram[4058]  = 72;
  ram[4059]  = 72;
  ram[4060]  = 72;
  ram[4061]  = 72;
  ram[4062]  = 72;
  ram[4063]  = 72;
  ram[4064]  = 72;
  ram[4065]  = 72;
  ram[4066]  = 72;
  ram[4067]  = 72;
  ram[4068]  = 71;
  ram[4069]  = 71;
  ram[4070]  = 72;
  ram[4071]  = 72;
  ram[4072]  = 72;
  ram[4073]  = 72;
  ram[4074]  = 72;
  ram[4075]  = 72;
  ram[4076]  = 72;
  ram[4077]  = 72;
  ram[4078]  = 73;
  ram[4079]  = 73;
  ram[4080]  = 73;
  ram[4081]  = 73;
  ram[4082]  = 72;
  ram[4083]  = 72;
  ram[4084]  = 72;
  ram[4085]  = 73;
  ram[4086]  = 73;
  ram[4087]  = 73;
  ram[4088]  = 73;
  ram[4089]  = 73;
  ram[4090]  = 72;
  ram[4091]  = 72;
  ram[4092]  = 71;
  ram[4093]  = 71;
  ram[4094]  = 70;
  ram[4095]  = 69;
end

always @(posedge clock) begin
  dout <= ram[address];
end

endmodule
