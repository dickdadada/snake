module rom_snakeb (clock, address, q);
input clock;
output [7:0] q;
input [11:0] address;
reg [7:0] dout;
reg [7:0] ram [4095:0];
assign q = dout;

initial begin
  ram[0]  = 72;
  ram[1]  = 77;
  ram[2]  = 78;
  ram[3]  = 78;
  ram[4]  = 80;
  ram[5]  = 78;
  ram[6]  = 80;
  ram[7]  = 80;
  ram[8]  = 77;
  ram[9]  = 77;
  ram[10]  = 77;
  ram[11]  = 77;
  ram[12]  = 77;
  ram[13]  = 77;
  ram[14]  = 79;
  ram[15]  = 79;
  ram[16]  = 78;
  ram[17]  = 78;
  ram[18]  = 78;
  ram[19]  = 78;
  ram[20]  = 80;
  ram[21]  = 80;
  ram[22]  = 80;
  ram[23]  = 80;
  ram[24]  = 80;
  ram[25]  = 80;
  ram[26]  = 78;
  ram[27]  = 78;
  ram[28]  = 78;
  ram[29]  = 78;
  ram[30]  = 76;
  ram[31]  = 76;
  ram[32]  = 78;
  ram[33]  = 78;
  ram[34]  = 78;
  ram[35]  = 78;
  ram[36]  = 78;
  ram[37]  = 78;
  ram[38]  = 78;
  ram[39]  = 78;
  ram[40]  = 78;
  ram[41]  = 78;
  ram[42]  = 78;
  ram[43]  = 78;
  ram[44]  = 78;
  ram[45]  = 78;
  ram[46]  = 78;
  ram[47]  = 78;
  ram[48]  = 76;
  ram[49]  = 76;
  ram[50]  = 78;
  ram[51]  = 78;
  ram[52]  = 78;
  ram[53]  = 78;
  ram[54]  = 78;
  ram[55]  = 78;
  ram[56]  = 77;
  ram[57]  = 78;
  ram[58]  = 78;
  ram[59]  = 78;
  ram[60]  = 78;
  ram[61]  = 78;
  ram[62]  = 75;
  ram[63]  = 73;
  ram[64]  = 75;
  ram[65]  = 79;
  ram[66]  = 80;
  ram[67]  = 80;
  ram[68]  = 83;
  ram[69]  = 81;
  ram[70]  = 83;
  ram[71]  = 82;
  ram[72]  = 80;
  ram[73]  = 80;
  ram[74]  = 80;
  ram[75]  = 80;
  ram[76]  = 80;
  ram[77]  = 80;
  ram[78]  = 82;
  ram[79]  = 82;
  ram[80]  = 80;
  ram[81]  = 80;
  ram[82]  = 80;
  ram[83]  = 80;
  ram[84]  = 82;
  ram[85]  = 82;
  ram[86]  = 82;
  ram[87]  = 82;
  ram[88]  = 82;
  ram[89]  = 82;
  ram[90]  = 80;
  ram[91]  = 80;
  ram[92]  = 80;
  ram[93]  = 80;
  ram[94]  = 78;
  ram[95]  = 78;
  ram[96]  = 80;
  ram[97]  = 80;
  ram[98]  = 80;
  ram[99]  = 80;
  ram[100]  = 80;
  ram[101]  = 80;
  ram[102]  = 80;
  ram[103]  = 80;
  ram[104]  = 80;
  ram[105]  = 80;
  ram[106]  = 80;
  ram[107]  = 80;
  ram[108]  = 80;
  ram[109]  = 80;
  ram[110]  = 80;
  ram[111]  = 80;
  ram[112]  = 78;
  ram[113]  = 78;
  ram[114]  = 80;
  ram[115]  = 80;
  ram[116]  = 80;
  ram[117]  = 80;
  ram[118]  = 80;
  ram[119]  = 80;
  ram[120]  = 80;
  ram[121]  = 80;
  ram[122]  = 80;
  ram[123]  = 80;
  ram[124]  = 81;
  ram[125]  = 81;
  ram[126]  = 78;
  ram[127]  = 75;
  ram[128]  = 76;
  ram[129]  = 80;
  ram[130]  = 80;
  ram[131]  = 81;
  ram[132]  = 84;
  ram[133]  = 83;
  ram[134]  = 83;
  ram[135]  = 83;
  ram[136]  = 82;
  ram[137]  = 82;
  ram[138]  = 81;
  ram[139]  = 81;
  ram[140]  = 81;
  ram[141]  = 81;
  ram[142]  = 83;
  ram[143]  = 83;
  ram[144]  = 81;
  ram[145]  = 81;
  ram[146]  = 81;
  ram[147]  = 81;
  ram[148]  = 83;
  ram[149]  = 83;
  ram[150]  = 83;
  ram[151]  = 83;
  ram[152]  = 83;
  ram[153]  = 83;
  ram[154]  = 83;
  ram[155]  = 83;
  ram[156]  = 81;
  ram[157]  = 81;
  ram[158]  = 81;
  ram[159]  = 81;
  ram[160]  = 81;
  ram[161]  = 81;
  ram[162]  = 81;
  ram[163]  = 81;
  ram[164]  = 81;
  ram[165]  = 81;
  ram[166]  = 81;
  ram[167]  = 81;
  ram[168]  = 81;
  ram[169]  = 81;
  ram[170]  = 81;
  ram[171]  = 81;
  ram[172]  = 81;
  ram[173]  = 81;
  ram[174]  = 81;
  ram[175]  = 81;
  ram[176]  = 79;
  ram[177]  = 79;
  ram[178]  = 81;
  ram[179]  = 81;
  ram[180]  = 81;
  ram[181]  = 81;
  ram[182]  = 81;
  ram[183]  = 81;
  ram[184]  = 81;
  ram[185]  = 81;
  ram[186]  = 81;
  ram[187]  = 81;
  ram[188]  = 81;
  ram[189]  = 82;
  ram[190]  = 78;
  ram[191]  = 76;
  ram[192]  = 76;
  ram[193]  = 79;
  ram[194]  = 79;
  ram[195]  = 80;
  ram[196]  = 84;
  ram[197]  = 83;
  ram[198]  = 83;
  ram[199]  = 82;
  ram[200]  = 82;
  ram[201]  = 82;
  ram[202]  = 82;
  ram[203]  = 82;
  ram[204]  = 82;
  ram[205]  = 82;
  ram[206]  = 84;
  ram[207]  = 84;
  ram[208]  = 81;
  ram[209]  = 81;
  ram[210]  = 81;
  ram[211]  = 81;
  ram[212]  = 83;
  ram[213]  = 83;
  ram[214]  = 83;
  ram[215]  = 83;
  ram[216]  = 83;
  ram[217]  = 83;
  ram[218]  = 83;
  ram[219]  = 83;
  ram[220]  = 81;
  ram[221]  = 81;
  ram[222]  = 81;
  ram[223]  = 81;
  ram[224]  = 81;
  ram[225]  = 81;
  ram[226]  = 81;
  ram[227]  = 81;
  ram[228]  = 81;
  ram[229]  = 81;
  ram[230]  = 81;
  ram[231]  = 81;
  ram[232]  = 81;
  ram[233]  = 81;
  ram[234]  = 81;
  ram[235]  = 81;
  ram[236]  = 81;
  ram[237]  = 81;
  ram[238]  = 81;
  ram[239]  = 81;
  ram[240]  = 79;
  ram[241]  = 79;
  ram[242]  = 81;
  ram[243]  = 81;
  ram[244]  = 81;
  ram[245]  = 81;
  ram[246]  = 81;
  ram[247]  = 81;
  ram[248]  = 80;
  ram[249]  = 81;
  ram[250]  = 81;
  ram[251]  = 80;
  ram[252]  = 81;
  ram[253]  = 81;
  ram[254]  = 78;
  ram[255]  = 76;
  ram[256]  = 76;
  ram[257]  = 80;
  ram[258]  = 80;
  ram[259]  = 80;
  ram[260]  = 84;
  ram[261]  = 83;
  ram[262]  = 83;
  ram[263]  = 82;
  ram[264]  = 82;
  ram[265]  = 82;
  ram[266]  = 82;
  ram[267]  = 82;
  ram[268]  = 82;
  ram[269]  = 82;
  ram[270]  = 84;
  ram[271]  = 84;
  ram[272]  = 82;
  ram[273]  = 82;
  ram[274]  = 82;
  ram[275]  = 82;
  ram[276]  = 84;
  ram[277]  = 84;
  ram[278]  = 84;
  ram[279]  = 84;
  ram[280]  = 84;
  ram[281]  = 84;
  ram[282]  = 84;
  ram[283]  = 84;
  ram[284]  = 82;
  ram[285]  = 82;
  ram[286]  = 82;
  ram[287]  = 82;
  ram[288]  = 82;
  ram[289]  = 82;
  ram[290]  = 82;
  ram[291]  = 82;
  ram[292]  = 82;
  ram[293]  = 82;
  ram[294]  = 82;
  ram[295]  = 82;
  ram[296]  = 82;
  ram[297]  = 82;
  ram[298]  = 82;
  ram[299]  = 82;
  ram[300]  = 82;
  ram[301]  = 82;
  ram[302]  = 82;
  ram[303]  = 82;
  ram[304]  = 82;
  ram[305]  = 82;
  ram[306]  = 82;
  ram[307]  = 82;
  ram[308]  = 82;
  ram[309]  = 82;
  ram[310]  = 84;
  ram[311]  = 84;
  ram[312]  = 83;
  ram[313]  = 83;
  ram[314]  = 81;
  ram[315]  = 81;
  ram[316]  = 81;
  ram[317]  = 82;
  ram[318]  = 80;
  ram[319]  = 78;
  ram[320]  = 76;
  ram[321]  = 80;
  ram[322]  = 80;
  ram[323]  = 80;
  ram[324]  = 84;
  ram[325]  = 82;
  ram[326]  = 83;
  ram[327]  = 82;
  ram[328]  = 81;
  ram[329]  = 81;
  ram[330]  = 81;
  ram[331]  = 81;
  ram[332]  = 80;
  ram[333]  = 81;
  ram[334]  = 83;
  ram[335]  = 83;
  ram[336]  = 81;
  ram[337]  = 81;
  ram[338]  = 81;
  ram[339]  = 81;
  ram[340]  = 83;
  ram[341]  = 83;
  ram[342]  = 83;
  ram[343]  = 83;
  ram[344]  = 83;
  ram[345]  = 83;
  ram[346]  = 83;
  ram[347]  = 83;
  ram[348]  = 81;
  ram[349]  = 81;
  ram[350]  = 81;
  ram[351]  = 81;
  ram[352]  = 81;
  ram[353]  = 81;
  ram[354]  = 81;
  ram[355]  = 81;
  ram[356]  = 81;
  ram[357]  = 81;
  ram[358]  = 81;
  ram[359]  = 81;
  ram[360]  = 81;
  ram[361]  = 81;
  ram[362]  = 81;
  ram[363]  = 81;
  ram[364]  = 81;
  ram[365]  = 81;
  ram[366]  = 81;
  ram[367]  = 81;
  ram[368]  = 81;
  ram[369]  = 81;
  ram[370]  = 81;
  ram[371]  = 81;
  ram[372]  = 81;
  ram[373]  = 81;
  ram[374]  = 83;
  ram[375]  = 83;
  ram[376]  = 83;
  ram[377]  = 83;
  ram[378]  = 81;
  ram[379]  = 81;
  ram[380]  = 81;
  ram[381]  = 81;
  ram[382]  = 80;
  ram[383]  = 78;
  ram[384]  = 75;
  ram[385]  = 79;
  ram[386]  = 80;
  ram[387]  = 80;
  ram[388]  = 83;
  ram[389]  = 82;
  ram[390]  = 83;
  ram[391]  = 82;
  ram[392]  = 80;
  ram[393]  = 80;
  ram[394]  = 80;
  ram[395]  = 80;
  ram[396]  = 82;
  ram[397]  = 82;
  ram[398]  = 84;
  ram[399]  = 82;
  ram[400]  = 80;
  ram[401]  = 80;
  ram[402]  = 80;
  ram[403]  = 80;
  ram[404]  = 82;
  ram[405]  = 82;
  ram[406]  = 82;
  ram[407]  = 82;
  ram[408]  = 82;
  ram[409]  = 82;
  ram[410]  = 82;
  ram[411]  = 82;
  ram[412]  = 82;
  ram[413]  = 82;
  ram[414]  = 82;
  ram[415]  = 82;
  ram[416]  = 82;
  ram[417]  = 82;
  ram[418]  = 82;
  ram[419]  = 82;
  ram[420]  = 82;
  ram[421]  = 82;
  ram[422]  = 82;
  ram[423]  = 82;
  ram[424]  = 82;
  ram[425]  = 82;
  ram[426]  = 82;
  ram[427]  = 82;
  ram[428]  = 80;
  ram[429]  = 80;
  ram[430]  = 80;
  ram[431]  = 80;
  ram[432]  = 80;
  ram[433]  = 80;
  ram[434]  = 80;
  ram[435]  = 80;
  ram[436]  = 82;
  ram[437]  = 82;
  ram[438]  = 82;
  ram[439]  = 82;
  ram[440]  = 83;
  ram[441]  = 83;
  ram[442]  = 83;
  ram[443]  = 82;
  ram[444]  = 81;
  ram[445]  = 81;
  ram[446]  = 79;
  ram[447]  = 77;
  ram[448]  = 75;
  ram[449]  = 80;
  ram[450]  = 81;
  ram[451]  = 81;
  ram[452]  = 84;
  ram[453]  = 82;
  ram[454]  = 83;
  ram[455]  = 84;
  ram[456]  = 84;
  ram[457]  = 82;
  ram[458]  = 81;
  ram[459]  = 81;
  ram[460]  = 83;
  ram[461]  = 83;
  ram[462]  = 85;
  ram[463]  = 83;
  ram[464]  = 83;
  ram[465]  = 81;
  ram[466]  = 81;
  ram[467]  = 81;
  ram[468]  = 83;
  ram[469]  = 83;
  ram[470]  = 83;
  ram[471]  = 83;
  ram[472]  = 83;
  ram[473]  = 83;
  ram[474]  = 83;
  ram[475]  = 83;
  ram[476]  = 83;
  ram[477]  = 83;
  ram[478]  = 83;
  ram[479]  = 83;
  ram[480]  = 83;
  ram[481]  = 83;
  ram[482]  = 83;
  ram[483]  = 83;
  ram[484]  = 83;
  ram[485]  = 83;
  ram[486]  = 83;
  ram[487]  = 83;
  ram[488]  = 83;
  ram[489]  = 83;
  ram[490]  = 83;
  ram[491]  = 83;
  ram[492]  = 81;
  ram[493]  = 81;
  ram[494]  = 81;
  ram[495]  = 81;
  ram[496]  = 81;
  ram[497]  = 81;
  ram[498]  = 81;
  ram[499]  = 81;
  ram[500]  = 83;
  ram[501]  = 83;
  ram[502]  = 83;
  ram[503]  = 83;
  ram[504]  = 83;
  ram[505]  = 84;
  ram[506]  = 84;
  ram[507]  = 83;
  ram[508]  = 81;
  ram[509]  = 82;
  ram[510]  = 80;
  ram[511]  = 78;
  ram[512]  = 75;
  ram[513]  = 78;
  ram[514]  = 80;
  ram[515]  = 79;
  ram[516]  = 82;
  ram[517]  = 82;
  ram[518]  = 84;
  ram[519]  = 82;
  ram[520]  = 82;
  ram[521]  = 82;
  ram[522]  = 80;
  ram[523]  = 80;
  ram[524]  = 82;
  ram[525]  = 82;
  ram[526]  = 84;
  ram[527]  = 82;
  ram[528]  = 82;
  ram[529]  = 80;
  ram[530]  = 81;
  ram[531]  = 81;
  ram[532]  = 80;
  ram[533]  = 80;
  ram[534]  = 82;
  ram[535]  = 83;
  ram[536]  = 82;
  ram[537]  = 82;
  ram[538]  = 82;
  ram[539]  = 82;
  ram[540]  = 82;
  ram[541]  = 82;
  ram[542]  = 82;
  ram[543]  = 82;
  ram[544]  = 82;
  ram[545]  = 82;
  ram[546]  = 82;
  ram[547]  = 82;
  ram[548]  = 82;
  ram[549]  = 82;
  ram[550]  = 82;
  ram[551]  = 82;
  ram[552]  = 81;
  ram[553]  = 82;
  ram[554]  = 82;
  ram[555]  = 82;
  ram[556]  = 80;
  ram[557]  = 80;
  ram[558]  = 80;
  ram[559]  = 80;
  ram[560]  = 80;
  ram[561]  = 80;
  ram[562]  = 80;
  ram[563]  = 80;
  ram[564]  = 82;
  ram[565]  = 82;
  ram[566]  = 82;
  ram[567]  = 81;
  ram[568]  = 81;
  ram[569]  = 82;
  ram[570]  = 82;
  ram[571]  = 82;
  ram[572]  = 80;
  ram[573]  = 81;
  ram[574]  = 79;
  ram[575]  = 78;
  ram[576]  = 76;
  ram[577]  = 80;
  ram[578]  = 82;
  ram[579]  = 81;
  ram[580]  = 84;
  ram[581]  = 84;
  ram[582]  = 85;
  ram[583]  = 85;
  ram[584]  = 83;
  ram[585]  = 83;
  ram[586]  = 81;
  ram[587]  = 81;
  ram[588]  = 83;
  ram[589]  = 83;
  ram[590]  = 85;
  ram[591]  = 85;
  ram[592]  = 83;
  ram[593]  = 82;
  ram[594]  = 82;
  ram[595]  = 82;
  ram[596]  = 81;
  ram[597]  = 81;
  ram[598]  = 83;
  ram[599]  = 83;
  ram[600]  = 84;
  ram[601]  = 84;
  ram[602]  = 84;
  ram[603]  = 84;
  ram[604]  = 84;
  ram[605]  = 84;
  ram[606]  = 84;
  ram[607]  = 83;
  ram[608]  = 84;
  ram[609]  = 84;
  ram[610]  = 84;
  ram[611]  = 84;
  ram[612]  = 84;
  ram[613]  = 85;
  ram[614]  = 85;
  ram[615]  = 85;
  ram[616]  = 85;
  ram[617]  = 85;
  ram[618]  = 85;
  ram[619]  = 85;
  ram[620]  = 83;
  ram[621]  = 83;
  ram[622]  = 83;
  ram[623]  = 83;
  ram[624]  = 82;
  ram[625]  = 82;
  ram[626]  = 82;
  ram[627]  = 82;
  ram[628]  = 84;
  ram[629]  = 84;
  ram[630]  = 84;
  ram[631]  = 83;
  ram[632]  = 83;
  ram[633]  = 84;
  ram[634]  = 84;
  ram[635]  = 83;
  ram[636]  = 81;
  ram[637]  = 81;
  ram[638]  = 80;
  ram[639]  = 78;
  ram[640]  = 78;
  ram[641]  = 81;
  ram[642]  = 82;
  ram[643]  = 81;
  ram[644]  = 84;
  ram[645]  = 86;
  ram[646]  = 85;
  ram[647]  = 85;
  ram[648]  = 83;
  ram[649]  = 83;
  ram[650]  = 81;
  ram[651]  = 81;
  ram[652]  = 83;
  ram[653]  = 83;
  ram[654]  = 85;
  ram[655]  = 85;
  ram[656]  = 84;
  ram[657]  = 84;
  ram[658]  = 81;
  ram[659]  = 81;
  ram[660]  = 81;
  ram[661]  = 81;
  ram[662]  = 81;
  ram[663]  = 81;
  ram[664]  = 83;
  ram[665]  = 83;
  ram[666]  = 83;
  ram[667]  = 83;
  ram[668]  = 85;
  ram[669]  = 85;
  ram[670]  = 85;
  ram[671]  = 85;
  ram[672]  = 85;
  ram[673]  = 85;
  ram[674]  = 85;
  ram[675]  = 84;
  ram[676]  = 84;
  ram[677]  = 84;
  ram[678]  = 82;
  ram[679]  = 82;
  ram[680]  = 82;
  ram[681]  = 82;
  ram[682]  = 82;
  ram[683]  = 82;
  ram[684]  = 82;
  ram[685]  = 82;
  ram[686]  = 80;
  ram[687]  = 80;
  ram[688]  = 81;
  ram[689]  = 81;
  ram[690]  = 83;
  ram[691]  = 84;
  ram[692]  = 83;
  ram[693]  = 83;
  ram[694]  = 83;
  ram[695]  = 83;
  ram[696]  = 83;
  ram[697]  = 84;
  ram[698]  = 84;
  ram[699]  = 83;
  ram[700]  = 83;
  ram[701]  = 83;
  ram[702]  = 80;
  ram[703]  = 78;
  ram[704]  = 77;
  ram[705]  = 80;
  ram[706]  = 81;
  ram[707]  = 80;
  ram[708]  = 85;
  ram[709]  = 85;
  ram[710]  = 83;
  ram[711]  = 84;
  ram[712]  = 82;
  ram[713]  = 82;
  ram[714]  = 80;
  ram[715]  = 80;
  ram[716]  = 82;
  ram[717]  = 82;
  ram[718]  = 84;
  ram[719]  = 84;
  ram[720]  = 83;
  ram[721]  = 83;
  ram[722]  = 80;
  ram[723]  = 80;
  ram[724]  = 80;
  ram[725]  = 80;
  ram[726]  = 80;
  ram[727]  = 79;
  ram[728]  = 80;
  ram[729]  = 81;
  ram[730]  = 81;
  ram[731]  = 81;
  ram[732]  = 83;
  ram[733]  = 84;
  ram[734]  = 84;
  ram[735]  = 84;
  ram[736]  = 87;
  ram[737]  = 87;
  ram[738]  = 87;
  ram[739]  = 86;
  ram[740]  = 86;
  ram[741]  = 86;
  ram[742]  = 84;
  ram[743]  = 84;
  ram[744]  = 83;
  ram[745]  = 83;
  ram[746]  = 83;
  ram[747]  = 83;
  ram[748]  = 84;
  ram[749]  = 84;
  ram[750]  = 82;
  ram[751]  = 82;
  ram[752]  = 80;
  ram[753]  = 80;
  ram[754]  = 82;
  ram[755]  = 82;
  ram[756]  = 82;
  ram[757]  = 82;
  ram[758]  = 82;
  ram[759]  = 82;
  ram[760]  = 81;
  ram[761]  = 82;
  ram[762]  = 82;
  ram[763]  = 82;
  ram[764]  = 82;
  ram[765]  = 82;
  ram[766]  = 79;
  ram[767]  = 78;
  ram[768]  = 77;
  ram[769]  = 79;
  ram[770]  = 81;
  ram[771]  = 79;
  ram[772]  = 84;
  ram[773]  = 84;
  ram[774]  = 83;
  ram[775]  = 84;
  ram[776]  = 82;
  ram[777]  = 82;
  ram[778]  = 80;
  ram[779]  = 80;
  ram[780]  = 82;
  ram[781]  = 82;
  ram[782]  = 84;
  ram[783]  = 84;
  ram[784]  = 83;
  ram[785]  = 82;
  ram[786]  = 79;
  ram[787]  = 79;
  ram[788]  = 80;
  ram[789]  = 80;
  ram[790]  = 79;
  ram[791]  = 78;
  ram[792]  = 81;
  ram[793]  = 81;
  ram[794]  = 81;
  ram[795]  = 82;
  ram[796]  = 84;
  ram[797]  = 84;
  ram[798]  = 86;
  ram[799]  = 86;
  ram[800]  = 82;
  ram[801]  = 83;
  ram[802]  = 83;
  ram[803]  = 83;
  ram[804]  = 83;
  ram[805]  = 83;
  ram[806]  = 83;
  ram[807]  = 83;
  ram[808]  = 81;
  ram[809]  = 81;
  ram[810]  = 81;
  ram[811]  = 81;
  ram[812]  = 81;
  ram[813]  = 81;
  ram[814]  = 79;
  ram[815]  = 79;
  ram[816]  = 82;
  ram[817]  = 83;
  ram[818]  = 83;
  ram[819]  = 83;
  ram[820]  = 83;
  ram[821]  = 83;
  ram[822]  = 85;
  ram[823]  = 85;
  ram[824]  = 83;
  ram[825]  = 84;
  ram[826]  = 82;
  ram[827]  = 81;
  ram[828]  = 81;
  ram[829]  = 82;
  ram[830]  = 81;
  ram[831]  = 80;
  ram[832]  = 77;
  ram[833]  = 79;
  ram[834]  = 81;
  ram[835]  = 80;
  ram[836]  = 85;
  ram[837]  = 85;
  ram[838]  = 84;
  ram[839]  = 84;
  ram[840]  = 82;
  ram[841]  = 82;
  ram[842]  = 80;
  ram[843]  = 80;
  ram[844]  = 82;
  ram[845]  = 82;
  ram[846]  = 84;
  ram[847]  = 84;
  ram[848]  = 82;
  ram[849]  = 82;
  ram[850]  = 80;
  ram[851]  = 80;
  ram[852]  = 80;
  ram[853]  = 80;
  ram[854]  = 80;
  ram[855]  = 80;
  ram[856]  = 83;
  ram[857]  = 83;
  ram[858]  = 82;
  ram[859]  = 82;
  ram[860]  = 84;
  ram[861]  = 84;
  ram[862]  = 85;
  ram[863]  = 85;
  ram[864]  = 85;
  ram[865]  = 85;
  ram[866]  = 85;
  ram[867]  = 86;
  ram[868]  = 86;
  ram[869]  = 87;
  ram[870]  = 87;
  ram[871]  = 88;
  ram[872]  = 85;
  ram[873]  = 85;
  ram[874]  = 85;
  ram[875]  = 85;
  ram[876]  = 85;
  ram[877]  = 85;
  ram[878]  = 83;
  ram[879]  = 83;
  ram[880]  = 83;
  ram[881]  = 83;
  ram[882]  = 83;
  ram[883]  = 83;
  ram[884]  = 83;
  ram[885]  = 83;
  ram[886]  = 85;
  ram[887]  = 85;
  ram[888]  = 85;
  ram[889]  = 85;
  ram[890]  = 83;
  ram[891]  = 82;
  ram[892]  = 81;
  ram[893]  = 81;
  ram[894]  = 81;
  ram[895]  = 79;
  ram[896]  = 75;
  ram[897]  = 78;
  ram[898]  = 80;
  ram[899]  = 79;
  ram[900]  = 84;
  ram[901]  = 84;
  ram[902]  = 83;
  ram[903]  = 84;
  ram[904]  = 82;
  ram[905]  = 82;
  ram[906]  = 80;
  ram[907]  = 80;
  ram[908]  = 81;
  ram[909]  = 81;
  ram[910]  = 83;
  ram[911]  = 83;
  ram[912]  = 81;
  ram[913]  = 81;
  ram[914]  = 79;
  ram[915]  = 79;
  ram[916]  = 79;
  ram[917]  = 79;
  ram[918]  = 79;
  ram[919]  = 80;
  ram[920]  = 81;
  ram[921]  = 81;
  ram[922]  = 81;
  ram[923]  = 81;
  ram[924]  = 83;
  ram[925]  = 83;
  ram[926]  = 85;
  ram[927]  = 85;
  ram[928]  = 85;
  ram[929]  = 85;
  ram[930]  = 83;
  ram[931]  = 83;
  ram[932]  = 83;
  ram[933]  = 83;
  ram[934]  = 83;
  ram[935]  = 83;
  ram[936]  = 81;
  ram[937]  = 81;
  ram[938]  = 81;
  ram[939]  = 81;
  ram[940]  = 81;
  ram[941]  = 81;
  ram[942]  = 79;
  ram[943]  = 79;
  ram[944]  = 82;
  ram[945]  = 82;
  ram[946]  = 82;
  ram[947]  = 82;
  ram[948]  = 82;
  ram[949]  = 82;
  ram[950]  = 84;
  ram[951]  = 84;
  ram[952]  = 84;
  ram[953]  = 85;
  ram[954]  = 82;
  ram[955]  = 81;
  ram[956]  = 81;
  ram[957]  = 81;
  ram[958]  = 80;
  ram[959]  = 79;
  ram[960]  = 75;
  ram[961]  = 76;
  ram[962]  = 76;
  ram[963]  = 77;
  ram[964]  = 82;
  ram[965]  = 83;
  ram[966]  = 80;
  ram[967]  = 79;
  ram[968]  = 75;
  ram[969]  = 73;
  ram[970]  = 73;
  ram[971]  = 75;
  ram[972]  = 76;
  ram[973]  = 78;
  ram[974]  = 82;
  ram[975]  = 82;
  ram[976]  = 75;
  ram[977]  = 76;
  ram[978]  = 80;
  ram[979]  = 80;
  ram[980]  = 80;
  ram[981]  = 78;
  ram[982]  = 80;
  ram[983]  = 79;
  ram[984]  = 77;
  ram[985]  = 78;
  ram[986]  = 80;
  ram[987]  = 80;
  ram[988]  = 79;
  ram[989]  = 80;
  ram[990]  = 80;
  ram[991]  = 80;
  ram[992]  = 81;
  ram[993]  = 81;
  ram[994]  = 80;
  ram[995]  = 79;
  ram[996]  = 80;
  ram[997]  = 80;
  ram[998]  = 77;
  ram[999]  = 77;
  ram[1000]  = 78;
  ram[1001]  = 78;
  ram[1002]  = 78;
  ram[1003]  = 80;
  ram[1004]  = 81;
  ram[1005]  = 81;
  ram[1006]  = 77;
  ram[1007]  = 77;
  ram[1008]  = 79;
  ram[1009]  = 79;
  ram[1010]  = 76;
  ram[1011]  = 75;
  ram[1012]  = 78;
  ram[1013]  = 80;
  ram[1014]  = 82;
  ram[1015]  = 82;
  ram[1016]  = 78;
  ram[1017]  = 76;
  ram[1018]  = 76;
  ram[1019]  = 77;
  ram[1020]  = 79;
  ram[1021]  = 82;
  ram[1022]  = 82;
  ram[1023]  = 80;
  ram[1024]  = 77;
  ram[1025]  = 77;
  ram[1026]  = 74;
  ram[1027]  = 72;
  ram[1028]  = 82;
  ram[1029]  = 79;
  ram[1030]  = 76;
  ram[1031]  = 49;
  ram[1032]  = 44;
  ram[1033]  = 46;
  ram[1034]  = 47;
  ram[1035]  = 46;
  ram[1036]  = 55;
  ram[1037]  = 54;
  ram[1038]  = 77;
  ram[1039]  = 77;
  ram[1040]  = 60;
  ram[1041]  = 52;
  ram[1042]  = 78;
  ram[1043]  = 81;
  ram[1044]  = 83;
  ram[1045]  = 77;
  ram[1046]  = 79;
  ram[1047]  = 73;
  ram[1048]  = 56;
  ram[1049]  = 64;
  ram[1050]  = 76;
  ram[1051]  = 80;
  ram[1052]  = 71;
  ram[1053]  = 60;
  ram[1054]  = 43;
  ram[1055]  = 50;
  ram[1056]  = 53;
  ram[1057]  = 52;
  ram[1058]  = 52;
  ram[1059]  = 68;
  ram[1060]  = 74;
  ram[1061]  = 72;
  ram[1062]  = 63;
  ram[1063]  = 52;
  ram[1064]  = 62;
  ram[1065]  = 72;
  ram[1066]  = 73;
  ram[1067]  = 75;
  ram[1068]  = 76;
  ram[1069]  = 77;
  ram[1070]  = 53;
  ram[1071]  = 50;
  ram[1072]  = 76;
  ram[1073]  = 71;
  ram[1074]  = 40;
  ram[1075]  = 48;
  ram[1076]  = 47;
  ram[1077]  = 58;
  ram[1078]  = 57;
  ram[1079]  = 58;
  ram[1080]  = 54;
  ram[1081]  = 55;
  ram[1082]  = 48;
  ram[1083]  = 63;
  ram[1084]  = 83;
  ram[1085]  = 83;
  ram[1086]  = 81;
  ram[1087]  = 81;
  ram[1088]  = 76;
  ram[1089]  = 79;
  ram[1090]  = 69;
  ram[1091]  = 72;
  ram[1092]  = 82;
  ram[1093]  = 65;
  ram[1094]  = 68;
  ram[1095]  = 124;
  ram[1096]  = 99;
  ram[1097]  = 97;
  ram[1098]  = 96;
  ram[1099]  = 113;
  ram[1100]  = 99;
  ram[1101]  = 137;
  ram[1102]  = 72;
  ram[1103]  = 47;
  ram[1104]  = 113;
  ram[1105]  = 121;
  ram[1106]  = 60;
  ram[1107]  = 85;
  ram[1108]  = 79;
  ram[1109]  = 81;
  ram[1110]  = 75;
  ram[1111]  = 82;
  ram[1112]  = 129;
  ram[1113]  = 90;
  ram[1114]  = 66;
  ram[1115]  = 75;
  ram[1116]  = 50;
  ram[1117]  = 97;
  ram[1118]  = 113;
  ram[1119]  = 101;
  ram[1120]  = 105;
  ram[1121]  = 110;
  ram[1122]  = 103;
  ram[1123]  = 55;
  ram[1124]  = 66;
  ram[1125]  = 59;
  ram[1126]  = 75;
  ram[1127]  = 128;
  ram[1128]  = 87;
  ram[1129]  = 61;
  ram[1130]  = 75;
  ram[1131]  = 70;
  ram[1132]  = 79;
  ram[1133]  = 60;
  ram[1134]  = 119;
  ram[1135]  = 133;
  ram[1136]  = 54;
  ram[1137]  = 56;
  ram[1138]  = 113;
  ram[1139]  = 86;
  ram[1140]  = 106;
  ram[1141]  = 101;
  ram[1142]  = 116;
  ram[1143]  = 108;
  ram[1144]  = 112;
  ram[1145]  = 104;
  ram[1146]  = 119;
  ram[1147]  = 78;
  ram[1148]  = 70;
  ram[1149]  = 82;
  ram[1150]  = 86;
  ram[1151]  = 83;
  ram[1152]  = 81;
  ram[1153]  = 72;
  ram[1154]  = 87;
  ram[1155]  = 75;
  ram[1156]  = 62;
  ram[1157]  = 36;
  ram[1158]  = 60;
  ram[1159]  = 175;
  ram[1160]  = 164;
  ram[1161]  = 169;
  ram[1162]  = 169;
  ram[1163]  = 169;
  ram[1164]  = 173;
  ram[1165]  = 179;
  ram[1166]  = 55;
  ram[1167]  = 6;
  ram[1168]  = 165;
  ram[1169]  = 169;
  ram[1170]  = 41;
  ram[1171]  = 73;
  ram[1172]  = 83;
  ram[1173]  = 74;
  ram[1174]  = 59;
  ram[1175]  = 86;
  ram[1176]  = 167;
  ram[1177]  = 106;
  ram[1178]  = 39;
  ram[1179]  = 47;
  ram[1180]  = 22;
  ram[1181]  = 141;
  ram[1182]  = 170;
  ram[1183]  = 165;
  ram[1184]  = 166;
  ram[1185]  = 166;
  ram[1186]  = 158;
  ram[1187]  = 20;
  ram[1188]  = 44;
  ram[1189]  = 54;
  ram[1190]  = 87;
  ram[1191]  = 179;
  ram[1192]  = 101;
  ram[1193]  = 50;
  ram[1194]  = 64;
  ram[1195]  = 78;
  ram[1196]  = 43;
  ram[1197]  = 7;
  ram[1198]  = 190;
  ram[1199]  = 194;
  ram[1200]  = 18;
  ram[1201]  = 36;
  ram[1202]  = 160;
  ram[1203]  = 138;
  ram[1204]  = 162;
  ram[1205]  = 163;
  ram[1206]  = 169;
  ram[1207]  = 166;
  ram[1208]  = 169;
  ram[1209]  = 171;
  ram[1210]  = 184;
  ram[1211]  = 88;
  ram[1212]  = 64;
  ram[1213]  = 80;
  ram[1214]  = 79;
  ram[1215]  = 75;
  ram[1216]  = 73;
  ram[1217]  = 80;
  ram[1218]  = 87;
  ram[1219]  = 73;
  ram[1220]  = 65;
  ram[1221]  = 139;
  ram[1222]  = 98;
  ram[1223]  = 55;
  ram[1224]  = 62;
  ram[1225]  = 64;
  ram[1226]  = 59;
  ram[1227]  = 67;
  ram[1228]  = 63;
  ram[1229]  = 79;
  ram[1230]  = 43;
  ram[1231]  = 9;
  ram[1232]  = 145;
  ram[1233]  = 152;
  ram[1234]  = 24;
  ram[1235]  = 62;
  ram[1236]  = 82;
  ram[1237]  = 80;
  ram[1238]  = 49;
  ram[1239]  = 68;
  ram[1240]  = 156;
  ram[1241]  = 71;
  ram[1242]  = 19;
  ram[1243]  = 104;
  ram[1244]  = 133;
  ram[1245]  = 60;
  ram[1246]  = 59;
  ram[1247]  = 62;
  ram[1248]  = 58;
  ram[1249]  = 52;
  ram[1250]  = 55;
  ram[1251]  = 141;
  ram[1252]  = 122;
  ram[1253]  = 33;
  ram[1254]  = 64;
  ram[1255]  = 161;
  ram[1256]  = 86;
  ram[1257]  = 45;
  ram[1258]  = 62;
  ram[1259]  = 49;
  ram[1260]  = 128;
  ram[1261]  = 147;
  ram[1262]  = 65;
  ram[1263]  = 78;
  ram[1264]  = 42;
  ram[1265]  = 35;
  ram[1266]  = 154;
  ram[1267]  = 99;
  ram[1268]  = 31;
  ram[1269]  = 47;
  ram[1270]  = 64;
  ram[1271]  = 54;
  ram[1272]  = 63;
  ram[1273]  = 66;
  ram[1274]  = 81;
  ram[1275]  = 59;
  ram[1276]  = 71;
  ram[1277]  = 75;
  ram[1278]  = 70;
  ram[1279]  = 75;
  ram[1280]  = 77;
  ram[1281]  = 82;
  ram[1282]  = 77;
  ram[1283]  = 67;
  ram[1284]  = 59;
  ram[1285]  = 173;
  ram[1286]  = 152;
  ram[1287]  = 17;
  ram[1288]  = 55;
  ram[1289]  = 63;
  ram[1290]  = 63;
  ram[1291]  = 52;
  ram[1292]  = 61;
  ram[1293]  = 57;
  ram[1294]  = 64;
  ram[1295]  = 23;
  ram[1296]  = 158;
  ram[1297]  = 153;
  ram[1298]  = 0;
  ram[1299]  = 28;
  ram[1300]  = 75;
  ram[1301]  = 73;
  ram[1302]  = 57;
  ram[1303]  = 71;
  ram[1304]  = 154;
  ram[1305]  = 86;
  ram[1306]  = 7;
  ram[1307]  = 122;
  ram[1308]  = 175;
  ram[1309]  = 58;
  ram[1310]  = 38;
  ram[1311]  = 55;
  ram[1312]  = 58;
  ram[1313]  = 37;
  ram[1314]  = 41;
  ram[1315]  = 162;
  ram[1316]  = 141;
  ram[1317]  = 15;
  ram[1318]  = 66;
  ram[1319]  = 165;
  ram[1320]  = 84;
  ram[1321]  = 40;
  ram[1322]  = 34;
  ram[1323]  = 0;
  ram[1324]  = 182;
  ram[1325]  = 196;
  ram[1326]  = 40;
  ram[1327]  = 56;
  ram[1328]  = 57;
  ram[1329]  = 39;
  ram[1330]  = 163;
  ram[1331]  = 121;
  ram[1332]  = 3;
  ram[1333]  = 38;
  ram[1334]  = 44;
  ram[1335]  = 48;
  ram[1336]  = 51;
  ram[1337]  = 54;
  ram[1338]  = 60;
  ram[1339]  = 67;
  ram[1340]  = 73;
  ram[1341]  = 72;
  ram[1342]  = 77;
  ram[1343]  = 73;
  ram[1344]  = 76;
  ram[1345]  = 82;
  ram[1346]  = 75;
  ram[1347]  = 65;
  ram[1348]  = 41;
  ram[1349]  = 168;
  ram[1350]  = 120;
  ram[1351]  = 38;
  ram[1352]  = 66;
  ram[1353]  = 76;
  ram[1354]  = 78;
  ram[1355]  = 73;
  ram[1356]  = 66;
  ram[1357]  = 82;
  ram[1358]  = 79;
  ram[1359]  = 28;
  ram[1360]  = 146;
  ram[1361]  = 125;
  ram[1362]  = 124;
  ram[1363]  = 150;
  ram[1364]  = 39;
  ram[1365]  = 59;
  ram[1366]  = 47;
  ram[1367]  = 74;
  ram[1368]  = 159;
  ram[1369]  = 67;
  ram[1370]  = 3;
  ram[1371]  = 103;
  ram[1372]  = 151;
  ram[1373]  = 53;
  ram[1374]  = 55;
  ram[1375]  = 73;
  ram[1376]  = 69;
  ram[1377]  = 55;
  ram[1378]  = 42;
  ram[1379]  = 146;
  ram[1380]  = 121;
  ram[1381]  = 6;
  ram[1382]  = 55;
  ram[1383]  = 157;
  ram[1384]  = 73;
  ram[1385]  = 21;
  ram[1386]  = 121;
  ram[1387]  = 172;
  ram[1388]  = 51;
  ram[1389]  = 58;
  ram[1390]  = 61;
  ram[1391]  = 68;
  ram[1392]  = 66;
  ram[1393]  = 24;
  ram[1394]  = 158;
  ram[1395]  = 117;
  ram[1396]  = 13;
  ram[1397]  = 63;
  ram[1398]  = 64;
  ram[1399]  = 63;
  ram[1400]  = 62;
  ram[1401]  = 69;
  ram[1402]  = 77;
  ram[1403]  = 79;
  ram[1404]  = 81;
  ram[1405]  = 72;
  ram[1406]  = 73;
  ram[1407]  = 70;
  ram[1408]  = 72;
  ram[1409]  = 76;
  ram[1410]  = 70;
  ram[1411]  = 61;
  ram[1412]  = 47;
  ram[1413]  = 161;
  ram[1414]  = 105;
  ram[1415]  = 0;
  ram[1416]  = 13;
  ram[1417]  = 19;
  ram[1418]  = 19;
  ram[1419]  = 30;
  ram[1420]  = 50;
  ram[1421]  = 68;
  ram[1422]  = 75;
  ram[1423]  = 30;
  ram[1424]  = 146;
  ram[1425]  = 130;
  ram[1426]  = 165;
  ram[1427]  = 175;
  ram[1428]  = 0;
  ram[1429]  = 34;
  ram[1430]  = 33;
  ram[1431]  = 73;
  ram[1432]  = 165;
  ram[1433]  = 80;
  ram[1434]  = 0;
  ram[1435]  = 102;
  ram[1436]  = 143;
  ram[1437]  = 12;
  ram[1438]  = 0;
  ram[1439]  = 17;
  ram[1440]  = 17;
  ram[1441]  = 0;
  ram[1442]  = 6;
  ram[1443]  = 143;
  ram[1444]  = 123;
  ram[1445]  = 4;
  ram[1446]  = 58;
  ram[1447]  = 164;
  ram[1448]  = 63;
  ram[1449]  = 0;
  ram[1450]  = 149;
  ram[1451]  = 204;
  ram[1452]  = 55;
  ram[1453]  = 51;
  ram[1454]  = 67;
  ram[1455]  = 77;
  ram[1456]  = 61;
  ram[1457]  = 39;
  ram[1458]  = 154;
  ram[1459]  = 100;
  ram[1460]  = 0;
  ram[1461]  = 17;
  ram[1462]  = 20;
  ram[1463]  = 22;
  ram[1464]  = 30;
  ram[1465]  = 51;
  ram[1466]  = 74;
  ram[1467]  = 80;
  ram[1468]  = 81;
  ram[1469]  = 78;
  ram[1470]  = 82;
  ram[1471]  = 80;
  ram[1472]  = 69;
  ram[1473]  = 68;
  ram[1474]  = 75;
  ram[1475]  = 57;
  ram[1476]  = 50;
  ram[1477]  = 153;
  ram[1478]  = 127;
  ram[1479]  = 150;
  ram[1480]  = 144;
  ram[1481]  = 165;
  ram[1482]  = 161;
  ram[1483]  = 183;
  ram[1484]  = 86;
  ram[1485]  = 52;
  ram[1486]  = 69;
  ram[1487]  = 21;
  ram[1488]  = 147;
  ram[1489]  = 143;
  ram[1490]  = 0;
  ram[1491]  = 6;
  ram[1492]  = 192;
  ram[1493]  = 160;
  ram[1494]  = 15;
  ram[1495]  = 60;
  ram[1496]  = 167;
  ram[1497]  = 77;
  ram[1498]  = 0;
  ram[1499]  = 94;
  ram[1500]  = 125;
  ram[1501]  = 120;
  ram[1502]  = 162;
  ram[1503]  = 163;
  ram[1504]  = 160;
  ram[1505]  = 156;
  ram[1506]  = 119;
  ram[1507]  = 129;
  ram[1508]  = 113;
  ram[1509]  = 0;
  ram[1510]  = 58;
  ram[1511]  = 140;
  ram[1512]  = 134;
  ram[1513]  = 186;
  ram[1514]  = 44;
  ram[1515]  = 21;
  ram[1516]  = 47;
  ram[1517]  = 67;
  ram[1518]  = 73;
  ram[1519]  = 65;
  ram[1520]  = 64;
  ram[1521]  = 32;
  ram[1522]  = 148;
  ram[1523]  = 108;
  ram[1524]  = 153;
  ram[1525]  = 155;
  ram[1526]  = 167;
  ram[1527]  = 169;
  ram[1528]  = 188;
  ram[1529]  = 108;
  ram[1530]  = 67;
  ram[1531]  = 84;
  ram[1532]  = 82;
  ram[1533]  = 76;
  ram[1534]  = 79;
  ram[1535]  = 73;
  ram[1536]  = 68;
  ram[1537]  = 72;
  ram[1538]  = 73;
  ram[1539]  = 66;
  ram[1540]  = 68;
  ram[1541]  = 182;
  ram[1542]  = 171;
  ram[1543]  = 169;
  ram[1544]  = 170;
  ram[1545]  = 177;
  ram[1546]  = 177;
  ram[1547]  = 193;
  ram[1548]  = 61;
  ram[1549]  = 16;
  ram[1550]  = 60;
  ram[1551]  = 19;
  ram[1552]  = 158;
  ram[1553]  = 160;
  ram[1554]  = 4;
  ram[1555]  = 50;
  ram[1556]  = 211;
  ram[1557]  = 162;
  ram[1558]  = 0;
  ram[1559]  = 42;
  ram[1560]  = 163;
  ram[1561]  = 93;
  ram[1562]  = 7;
  ram[1563]  = 104;
  ram[1564]  = 130;
  ram[1565]  = 137;
  ram[1566]  = 157;
  ram[1567]  = 174;
  ram[1568]  = 174;
  ram[1569]  = 167;
  ram[1570]  = 141;
  ram[1571]  = 134;
  ram[1572]  = 117;
  ram[1573]  = 3;
  ram[1574]  = 51;
  ram[1575]  = 137;
  ram[1576]  = 146;
  ram[1577]  = 183;
  ram[1578]  = 34;
  ram[1579]  = 0;
  ram[1580]  = 49;
  ram[1581]  = 69;
  ram[1582]  = 73;
  ram[1583]  = 77;
  ram[1584]  = 64;
  ram[1585]  = 35;
  ram[1586]  = 150;
  ram[1587]  = 120;
  ram[1588]  = 167;
  ram[1589]  = 174;
  ram[1590]  = 184;
  ram[1591]  = 182;
  ram[1592]  = 192;
  ram[1593]  = 102;
  ram[1594]  = 70;
  ram[1595]  = 81;
  ram[1596]  = 85;
  ram[1597]  = 84;
  ram[1598]  = 77;
  ram[1599]  = 78;
  ram[1600]  = 74;
  ram[1601]  = 69;
  ram[1602]  = 74;
  ram[1603]  = 70;
  ram[1604]  = 68;
  ram[1605]  = 30;
  ram[1606]  = 13;
  ram[1607]  = 16;
  ram[1608]  = 8;
  ram[1609]  = 19;
  ram[1610]  = 11;
  ram[1611]  = 0;
  ram[1612]  = 123;
  ram[1613]  = 201;
  ram[1614]  = 68;
  ram[1615]  = 3;
  ram[1616]  = 152;
  ram[1617]  = 166;
  ram[1618]  = 25;
  ram[1619]  = 57;
  ram[1620]  = 22;
  ram[1621]  = 46;
  ram[1622]  = 188;
  ram[1623]  = 153;
  ram[1624]  = 145;
  ram[1625]  = 86;
  ram[1626]  = 0;
  ram[1627]  = 106;
  ram[1628]  = 141;
  ram[1629]  = 7;
  ram[1630]  = 0;
  ram[1631]  = 6;
  ram[1632]  = 10;
  ram[1633]  = 2;
  ram[1634]  = 0;
  ram[1635]  = 138;
  ram[1636]  = 119;
  ram[1637]  = 1;
  ram[1638]  = 50;
  ram[1639]  = 157;
  ram[1640]  = 49;
  ram[1641]  = 0;
  ram[1642]  = 126;
  ram[1643]  = 199;
  ram[1644]  = 66;
  ram[1645]  = 48;
  ram[1646]  = 74;
  ram[1647]  = 75;
  ram[1648]  = 66;
  ram[1649]  = 34;
  ram[1650]  = 162;
  ram[1651]  = 99;
  ram[1652]  = 0;
  ram[1653]  = 10;
  ram[1654]  = 15;
  ram[1655]  = 19;
  ram[1656]  = 30;
  ram[1657]  = 56;
  ram[1658]  = 74;
  ram[1659]  = 81;
  ram[1660]  = 79;
  ram[1661]  = 76;
  ram[1662]  = 80;
  ram[1663]  = 75;
  ram[1664]  = 76;
  ram[1665]  = 78;
  ram[1666]  = 81;
  ram[1667]  = 77;
  ram[1668]  = 63;
  ram[1669]  = 65;
  ram[1670]  = 59;
  ram[1671]  = 59;
  ram[1672]  = 70;
  ram[1673]  = 68;
  ram[1674]  = 60;
  ram[1675]  = 31;
  ram[1676]  = 117;
  ram[1677]  = 180;
  ram[1678]  = 43;
  ram[1679]  = 0;
  ram[1680]  = 146;
  ram[1681]  = 153;
  ram[1682]  = 23;
  ram[1683]  = 57;
  ram[1684]  = 53;
  ram[1685]  = 75;
  ram[1686]  = 175;
  ram[1687]  = 140;
  ram[1688]  = 141;
  ram[1689]  = 72;
  ram[1690]  = 0;
  ram[1691]  = 109;
  ram[1692]  = 149;
  ram[1693]  = 37;
  ram[1694]  = 46;
  ram[1695]  = 64;
  ram[1696]  = 68;
  ram[1697]  = 46;
  ram[1698]  = 25;
  ram[1699]  = 156;
  ram[1700]  = 117;
  ram[1701]  = 0;
  ram[1702]  = 56;
  ram[1703]  = 162;
  ram[1704]  = 78;
  ram[1705]  = 0;
  ram[1706]  = 138;
  ram[1707]  = 182;
  ram[1708]  = 34;
  ram[1709]  = 35;
  ram[1710]  = 64;
  ram[1711]  = 69;
  ram[1712]  = 60;
  ram[1713]  = 40;
  ram[1714]  = 167;
  ram[1715]  = 126;
  ram[1716]  = 14;
  ram[1717]  = 52;
  ram[1718]  = 58;
  ram[1719]  = 64;
  ram[1720]  = 61;
  ram[1721]  = 69;
  ram[1722]  = 73;
  ram[1723]  = 80;
  ram[1724]  = 78;
  ram[1725]  = 77;
  ram[1726]  = 76;
  ram[1727]  = 76;
  ram[1728]  = 77;
  ram[1729]  = 84;
  ram[1730]  = 72;
  ram[1731]  = 75;
  ram[1732]  = 75;
  ram[1733]  = 63;
  ram[1734]  = 57;
  ram[1735]  = 53;
  ram[1736]  = 62;
  ram[1737]  = 52;
  ram[1738]  = 54;
  ram[1739]  = 19;
  ram[1740]  = 117;
  ram[1741]  = 178;
  ram[1742]  = 44;
  ram[1743]  = 0;
  ram[1744]  = 150;
  ram[1745]  = 158;
  ram[1746]  = 17;
  ram[1747]  = 59;
  ram[1748]  = 76;
  ram[1749]  = 54;
  ram[1750]  = 0;
  ram[1751]  = 36;
  ram[1752]  = 160;
  ram[1753]  = 79;
  ram[1754]  = 0;
  ram[1755]  = 103;
  ram[1756]  = 159;
  ram[1757]  = 46;
  ram[1758]  = 62;
  ram[1759]  = 80;
  ram[1760]  = 82;
  ram[1761]  = 55;
  ram[1762]  = 48;
  ram[1763]  = 149;
  ram[1764]  = 127;
  ram[1765]  = 0;
  ram[1766]  = 55;
  ram[1767]  = 169;
  ram[1768]  = 92;
  ram[1769]  = 39;
  ram[1770]  = 28;
  ram[1771]  = 0;
  ram[1772]  = 165;
  ram[1773]  = 200;
  ram[1774]  = 37;
  ram[1775]  = 51;
  ram[1776]  = 63;
  ram[1777]  = 33;
  ram[1778]  = 168;
  ram[1779]  = 127;
  ram[1780]  = 0;
  ram[1781]  = 50;
  ram[1782]  = 56;
  ram[1783]  = 55;
  ram[1784]  = 57;
  ram[1785]  = 56;
  ram[1786]  = 60;
  ram[1787]  = 72;
  ram[1788]  = 72;
  ram[1789]  = 76;
  ram[1790]  = 72;
  ram[1791]  = 73;
  ram[1792]  = 75;
  ram[1793]  = 70;
  ram[1794]  = 84;
  ram[1795]  = 71;
  ram[1796]  = 61;
  ram[1797]  = 64;
  ram[1798]  = 48;
  ram[1799]  = 52;
  ram[1800]  = 47;
  ram[1801]  = 46;
  ram[1802]  = 50;
  ram[1803]  = 40;
  ram[1804]  = 110;
  ram[1805]  = 179;
  ram[1806]  = 48;
  ram[1807]  = 0;
  ram[1808]  = 146;
  ram[1809]  = 156;
  ram[1810]  = 19;
  ram[1811]  = 65;
  ram[1812]  = 66;
  ram[1813]  = 76;
  ram[1814]  = 43;
  ram[1815]  = 69;
  ram[1816]  = 170;
  ram[1817]  = 77;
  ram[1818]  = 1;
  ram[1819]  = 108;
  ram[1820]  = 160;
  ram[1821]  = 57;
  ram[1822]  = 59;
  ram[1823]  = 81;
  ram[1824]  = 67;
  ram[1825]  = 57;
  ram[1826]  = 44;
  ram[1827]  = 162;
  ram[1828]  = 120;
  ram[1829]  = 0;
  ram[1830]  = 47;
  ram[1831]  = 168;
  ram[1832]  = 89;
  ram[1833]  = 47;
  ram[1834]  = 62;
  ram[1835]  = 43;
  ram[1836]  = 156;
  ram[1837]  = 170;
  ram[1838]  = 33;
  ram[1839]  = 64;
  ram[1840]  = 44;
  ram[1841]  = 26;
  ram[1842]  = 164;
  ram[1843]  = 100;
  ram[1844]  = 9;
  ram[1845]  = 33;
  ram[1846]  = 44;
  ram[1847]  = 38;
  ram[1848]  = 46;
  ram[1849]  = 55;
  ram[1850]  = 68;
  ram[1851]  = 56;
  ram[1852]  = 67;
  ram[1853]  = 70;
  ram[1854]  = 72;
  ram[1855]  = 73;
  ram[1856]  = 74;
  ram[1857]  = 73;
  ram[1858]  = 71;
  ram[1859]  = 69;
  ram[1860]  = 70;
  ram[1861]  = 197;
  ram[1862]  = 185;
  ram[1863]  = 176;
  ram[1864]  = 171;
  ram[1865]  = 176;
  ram[1866]  = 175;
  ram[1867]  = 197;
  ram[1868]  = 54;
  ram[1869]  = 7;
  ram[1870]  = 55;
  ram[1871]  = 10;
  ram[1872]  = 177;
  ram[1873]  = 172;
  ram[1874]  = 27;
  ram[1875]  = 69;
  ram[1876]  = 74;
  ram[1877]  = 69;
  ram[1878]  = 55;
  ram[1879]  = 91;
  ram[1880]  = 185;
  ram[1881]  = 105;
  ram[1882]  = 2;
  ram[1883]  = 127;
  ram[1884]  = 185;
  ram[1885]  = 70;
  ram[1886]  = 65;
  ram[1887]  = 81;
  ram[1888]  = 66;
  ram[1889]  = 59;
  ram[1890]  = 67;
  ram[1891]  = 181;
  ram[1892]  = 137;
  ram[1893]  = 0;
  ram[1894]  = 70;
  ram[1895]  = 182;
  ram[1896]  = 101;
  ram[1897]  = 52;
  ram[1898]  = 75;
  ram[1899]  = 75;
  ram[1900]  = 39;
  ram[1901]  = 0;
  ram[1902]  = 197;
  ram[1903]  = 205;
  ram[1904]  = 4;
  ram[1905]  = 38;
  ram[1906]  = 171;
  ram[1907]  = 137;
  ram[1908]  = 164;
  ram[1909]  = 170;
  ram[1910]  = 169;
  ram[1911]  = 173;
  ram[1912]  = 174;
  ram[1913]  = 178;
  ram[1914]  = 191;
  ram[1915]  = 85;
  ram[1916]  = 57;
  ram[1917]  = 69;
  ram[1918]  = 74;
  ram[1919]  = 69;
  ram[1920]  = 75;
  ram[1921]  = 75;
  ram[1922]  = 76;
  ram[1923]  = 61;
  ram[1924]  = 60;
  ram[1925]  = 149;
  ram[1926]  = 119;
  ram[1927]  = 137;
  ram[1928]  = 116;
  ram[1929]  = 131;
  ram[1930]  = 115;
  ram[1931]  = 148;
  ram[1932]  = 73;
  ram[1933]  = 54;
  ram[1934]  = 56;
  ram[1935]  = 43;
  ram[1936]  = 141;
  ram[1937]  = 152;
  ram[1938]  = 45;
  ram[1939]  = 62;
  ram[1940]  = 59;
  ram[1941]  = 67;
  ram[1942]  = 63;
  ram[1943]  = 87;
  ram[1944]  = 172;
  ram[1945]  = 81;
  ram[1946]  = 32;
  ram[1947]  = 107;
  ram[1948]  = 148;
  ram[1949]  = 63;
  ram[1950]  = 63;
  ram[1951]  = 71;
  ram[1952]  = 78;
  ram[1953]  = 64;
  ram[1954]  = 61;
  ram[1955]  = 150;
  ram[1956]  = 108;
  ram[1957]  = 26;
  ram[1958]  = 73;
  ram[1959]  = 163;
  ram[1960]  = 95;
  ram[1961]  = 61;
  ram[1962]  = 65;
  ram[1963]  = 73;
  ram[1964]  = 69;
  ram[1965]  = 41;
  ram[1966]  = 152;
  ram[1967]  = 169;
  ram[1968]  = 30;
  ram[1969]  = 43;
  ram[1970]  = 145;
  ram[1971]  = 97;
  ram[1972]  = 126;
  ram[1973]  = 118;
  ram[1974]  = 134;
  ram[1975]  = 120;
  ram[1976]  = 131;
  ram[1977]  = 114;
  ram[1978]  = 137;
  ram[1979]  = 71;
  ram[1980]  = 61;
  ram[1981]  = 72;
  ram[1982]  = 71;
  ram[1983]  = 73;
  ram[1984]  = 77;
  ram[1985]  = 76;
  ram[1986]  = 72;
  ram[1987]  = 70;
  ram[1988]  = 58;
  ram[1989]  = 37;
  ram[1990]  = 36;
  ram[1991]  = 30;
  ram[1992]  = 25;
  ram[1993]  = 21;
  ram[1994]  = 24;
  ram[1995]  = 32;
  ram[1996]  = 55;
  ram[1997]  = 70;
  ram[1998]  = 74;
  ram[1999]  = 65;
  ram[2000]  = 45;
  ram[2001]  = 39;
  ram[2002]  = 71;
  ram[2003]  = 68;
  ram[2004]  = 64;
  ram[2005]  = 62;
  ram[2006]  = 72;
  ram[2007]  = 58;
  ram[2008]  = 37;
  ram[2009]  = 54;
  ram[2010]  = 61;
  ram[2011]  = 39;
  ram[2012]  = 36;
  ram[2013]  = 53;
  ram[2014]  = 67;
  ram[2015]  = 75;
  ram[2016]  = 76;
  ram[2017]  = 73;
  ram[2018]  = 64;
  ram[2019]  = 32;
  ram[2020]  = 40;
  ram[2021]  = 55;
  ram[2022]  = 54;
  ram[2023]  = 44;
  ram[2024]  = 62;
  ram[2025]  = 74;
  ram[2026]  = 73;
  ram[2027]  = 74;
  ram[2028]  = 74;
  ram[2029]  = 70;
  ram[2030]  = 45;
  ram[2031]  = 41;
  ram[2032]  = 69;
  ram[2033]  = 57;
  ram[2034]  = 20;
  ram[2035]  = 23;
  ram[2036]  = 22;
  ram[2037]  = 26;
  ram[2038]  = 32;
  ram[2039]  = 32;
  ram[2040]  = 26;
  ram[2041]  = 26;
  ram[2042]  = 26;
  ram[2043]  = 42;
  ram[2044]  = 71;
  ram[2045]  = 73;
  ram[2046]  = 72;
  ram[2047]  = 72;
  ram[2048]  = 75;
  ram[2049]  = 75;
  ram[2050]  = 74;
  ram[2051]  = 71;
  ram[2052]  = 70;
  ram[2053]  = 70;
  ram[2054]  = 70;
  ram[2055]  = 70;
  ram[2056]  = 68;
  ram[2057]  = 70;
  ram[2058]  = 70;
  ram[2059]  = 71;
  ram[2060]  = 73;
  ram[2061]  = 75;
  ram[2062]  = 74;
  ram[2063]  = 71;
  ram[2064]  = 71;
  ram[2065]  = 72;
  ram[2066]  = 73;
  ram[2067]  = 71;
  ram[2068]  = 68;
  ram[2069]  = 68;
  ram[2070]  = 69;
  ram[2071]  = 69;
  ram[2072]  = 69;
  ram[2073]  = 69;
  ram[2074]  = 69;
  ram[2075]  = 68;
  ram[2076]  = 68;
  ram[2077]  = 68;
  ram[2078]  = 69;
  ram[2079]  = 74;
  ram[2080]  = 77;
  ram[2081]  = 77;
  ram[2082]  = 75;
  ram[2083]  = 74;
  ram[2084]  = 71;
  ram[2085]  = 69;
  ram[2086]  = 71;
  ram[2087]  = 73;
  ram[2088]  = 79;
  ram[2089]  = 77;
  ram[2090]  = 74;
  ram[2091]  = 72;
  ram[2092]  = 73;
  ram[2093]  = 76;
  ram[2094]  = 77;
  ram[2095]  = 77;
  ram[2096]  = 67;
  ram[2097]  = 66;
  ram[2098]  = 64;
  ram[2099]  = 66;
  ram[2100]  = 67;
  ram[2101]  = 68;
  ram[2102]  = 68;
  ram[2103]  = 69;
  ram[2104]  = 70;
  ram[2105]  = 70;
  ram[2106]  = 70;
  ram[2107]  = 72;
  ram[2108]  = 73;
  ram[2109]  = 74;
  ram[2110]  = 73;
  ram[2111]  = 73;
  ram[2112]  = 73;
  ram[2113]  = 73;
  ram[2114]  = 74;
  ram[2115]  = 74;
  ram[2116]  = 74;
  ram[2117]  = 74;
  ram[2118]  = 75;
  ram[2119]  = 76;
  ram[2120]  = 75;
  ram[2121]  = 76;
  ram[2122]  = 76;
  ram[2123]  = 74;
  ram[2124]  = 74;
  ram[2125]  = 75;
  ram[2126]  = 74;
  ram[2127]  = 74;
  ram[2128]  = 77;
  ram[2129]  = 78;
  ram[2130]  = 76;
  ram[2131]  = 76;
  ram[2132]  = 74;
  ram[2133]  = 72;
  ram[2134]  = 71;
  ram[2135]  = 71;
  ram[2136]  = 72;
  ram[2137]  = 72;
  ram[2138]  = 72;
  ram[2139]  = 72;
  ram[2140]  = 72;
  ram[2141]  = 72;
  ram[2142]  = 72;
  ram[2143]  = 72;
  ram[2144]  = 75;
  ram[2145]  = 74;
  ram[2146]  = 76;
  ram[2147]  = 76;
  ram[2148]  = 74;
  ram[2149]  = 71;
  ram[2150]  = 73;
  ram[2151]  = 75;
  ram[2152]  = 80;
  ram[2153]  = 80;
  ram[2154]  = 73;
  ram[2155]  = 71;
  ram[2156]  = 73;
  ram[2157]  = 75;
  ram[2158]  = 80;
  ram[2159]  = 80;
  ram[2160]  = 73;
  ram[2161]  = 73;
  ram[2162]  = 74;
  ram[2163]  = 74;
  ram[2164]  = 74;
  ram[2165]  = 74;
  ram[2166]  = 74;
  ram[2167]  = 74;
  ram[2168]  = 75;
  ram[2169]  = 76;
  ram[2170]  = 76;
  ram[2171]  = 76;
  ram[2172]  = 75;
  ram[2173]  = 74;
  ram[2174]  = 73;
  ram[2175]  = 73;
  ram[2176]  = 73;
  ram[2177]  = 73;
  ram[2178]  = 74;
  ram[2179]  = 74;
  ram[2180]  = 74;
  ram[2181]  = 74;
  ram[2182]  = 75;
  ram[2183]  = 75;
  ram[2184]  = 76;
  ram[2185]  = 76;
  ram[2186]  = 75;
  ram[2187]  = 73;
  ram[2188]  = 73;
  ram[2189]  = 74;
  ram[2190]  = 75;
  ram[2191]  = 75;
  ram[2192]  = 76;
  ram[2193]  = 77;
  ram[2194]  = 75;
  ram[2195]  = 75;
  ram[2196]  = 75;
  ram[2197]  = 75;
  ram[2198]  = 75;
  ram[2199]  = 75;
  ram[2200]  = 78;
  ram[2201]  = 78;
  ram[2202]  = 77;
  ram[2203]  = 77;
  ram[2204]  = 75;
  ram[2205]  = 75;
  ram[2206]  = 74;
  ram[2207]  = 74;
  ram[2208]  = 74;
  ram[2209]  = 73;
  ram[2210]  = 73;
  ram[2211]  = 73;
  ram[2212]  = 69;
  ram[2213]  = 68;
  ram[2214]  = 71;
  ram[2215]  = 75;
  ram[2216]  = 82;
  ram[2217]  = 82;
  ram[2218]  = 76;
  ram[2219]  = 71;
  ram[2220]  = 69;
  ram[2221]  = 69;
  ram[2222]  = 73;
  ram[2223]  = 75;
  ram[2224]  = 77;
  ram[2225]  = 75;
  ram[2226]  = 73;
  ram[2227]  = 73;
  ram[2228]  = 74;
  ram[2229]  = 74;
  ram[2230]  = 74;
  ram[2231]  = 73;
  ram[2232]  = 74;
  ram[2233]  = 75;
  ram[2234]  = 75;
  ram[2235]  = 75;
  ram[2236]  = 74;
  ram[2237]  = 73;
  ram[2238]  = 72;
  ram[2239]  = 72;
  ram[2240]  = 72;
  ram[2241]  = 72;
  ram[2242]  = 74;
  ram[2243]  = 74;
  ram[2244]  = 73;
  ram[2245]  = 73;
  ram[2246]  = 73;
  ram[2247]  = 73;
  ram[2248]  = 75;
  ram[2249]  = 74;
  ram[2250]  = 73;
  ram[2251]  = 72;
  ram[2252]  = 72;
  ram[2253]  = 73;
  ram[2254]  = 74;
  ram[2255]  = 74;
  ram[2256]  = 72;
  ram[2257]  = 72;
  ram[2258]  = 73;
  ram[2259]  = 72;
  ram[2260]  = 73;
  ram[2261]  = 73;
  ram[2262]  = 73;
  ram[2263]  = 75;
  ram[2264]  = 79;
  ram[2265]  = 79;
  ram[2266]  = 81;
  ram[2267]  = 79;
  ram[2268]  = 77;
  ram[2269]  = 74;
  ram[2270]  = 75;
  ram[2271]  = 74;
  ram[2272]  = 75;
  ram[2273]  = 72;
  ram[2274]  = 72;
  ram[2275]  = 70;
  ram[2276]  = 68;
  ram[2277]  = 67;
  ram[2278]  = 70;
  ram[2279]  = 75;
  ram[2280]  = 79;
  ram[2281]  = 79;
  ram[2282]  = 75;
  ram[2283]  = 70;
  ram[2284]  = 67;
  ram[2285]  = 64;
  ram[2286]  = 67;
  ram[2287]  = 70;
  ram[2288]  = 75;
  ram[2289]  = 73;
  ram[2290]  = 71;
  ram[2291]  = 71;
  ram[2292]  = 72;
  ram[2293]  = 73;
  ram[2294]  = 72;
  ram[2295]  = 72;
  ram[2296]  = 72;
  ram[2297]  = 73;
  ram[2298]  = 73;
  ram[2299]  = 73;
  ram[2300]  = 72;
  ram[2301]  = 71;
  ram[2302]  = 71;
  ram[2303]  = 70;
  ram[2304]  = 72;
  ram[2305]  = 72;
  ram[2306]  = 72;
  ram[2307]  = 72;
  ram[2308]  = 72;
  ram[2309]  = 71;
  ram[2310]  = 72;
  ram[2311]  = 71;
  ram[2312]  = 72;
  ram[2313]  = 72;
  ram[2314]  = 72;
  ram[2315]  = 72;
  ram[2316]  = 72;
  ram[2317]  = 71;
  ram[2318]  = 72;
  ram[2319]  = 71;
  ram[2320]  = 71;
  ram[2321]  = 69;
  ram[2322]  = 69;
  ram[2323]  = 69;
  ram[2324]  = 71;
  ram[2325]  = 71;
  ram[2326]  = 72;
  ram[2327]  = 74;
  ram[2328]  = 77;
  ram[2329]  = 76;
  ram[2330]  = 76;
  ram[2331]  = 76;
  ram[2332]  = 74;
  ram[2333]  = 72;
  ram[2334]  = 71;
  ram[2335]  = 71;
  ram[2336]  = 73;
  ram[2337]  = 72;
  ram[2338]  = 71;
  ram[2339]  = 70;
  ram[2340]  = 66;
  ram[2341]  = 64;
  ram[2342]  = 66;
  ram[2343]  = 70;
  ram[2344]  = 72;
  ram[2345]  = 72;
  ram[2346]  = 69;
  ram[2347]  = 65;
  ram[2348]  = 62;
  ram[2349]  = 62;
  ram[2350]  = 66;
  ram[2351]  = 70;
  ram[2352]  = 72;
  ram[2353]  = 71;
  ram[2354]  = 71;
  ram[2355]  = 71;
  ram[2356]  = 71;
  ram[2357]  = 71;
  ram[2358]  = 71;
  ram[2359]  = 71;
  ram[2360]  = 71;
  ram[2361]  = 71;
  ram[2362]  = 70;
  ram[2363]  = 70;
  ram[2364]  = 70;
  ram[2365]  = 69;
  ram[2366]  = 68;
  ram[2367]  = 67;
  ram[2368]  = 70;
  ram[2369]  = 70;
  ram[2370]  = 71;
  ram[2371]  = 71;
  ram[2372]  = 72;
  ram[2373]  = 71;
  ram[2374]  = 72;
  ram[2375]  = 71;
  ram[2376]  = 71;
  ram[2377]  = 71;
  ram[2378]  = 71;
  ram[2379]  = 72;
  ram[2380]  = 72;
  ram[2381]  = 71;
  ram[2382]  = 71;
  ram[2383]  = 71;
  ram[2384]  = 71;
  ram[2385]  = 71;
  ram[2386]  = 71;
  ram[2387]  = 71;
  ram[2388]  = 71;
  ram[2389]  = 71;
  ram[2390]  = 72;
  ram[2391]  = 74;
  ram[2392]  = 74;
  ram[2393]  = 74;
  ram[2394]  = 74;
  ram[2395]  = 74;
  ram[2396]  = 72;
  ram[2397]  = 70;
  ram[2398]  = 70;
  ram[2399]  = 70;
  ram[2400]  = 74;
  ram[2401]  = 73;
  ram[2402]  = 72;
  ram[2403]  = 71;
  ram[2404]  = 68;
  ram[2405]  = 65;
  ram[2406]  = 67;
  ram[2407]  = 70;
  ram[2408]  = 71;
  ram[2409]  = 71;
  ram[2410]  = 70;
  ram[2411]  = 67;
  ram[2412]  = 64;
  ram[2413]  = 64;
  ram[2414]  = 71;
  ram[2415]  = 74;
  ram[2416]  = 72;
  ram[2417]  = 71;
  ram[2418]  = 72;
  ram[2419]  = 72;
  ram[2420]  = 72;
  ram[2421]  = 71;
  ram[2422]  = 71;
  ram[2423]  = 71;
  ram[2424]  = 71;
  ram[2425]  = 71;
  ram[2426]  = 70;
  ram[2427]  = 70;
  ram[2428]  = 70;
  ram[2429]  = 69;
  ram[2430]  = 68;
  ram[2431]  = 68;
  ram[2432]  = 69;
  ram[2433]  = 70;
  ram[2434]  = 71;
  ram[2435]  = 71;
  ram[2436]  = 72;
  ram[2437]  = 71;
  ram[2438]  = 71;
  ram[2439]  = 70;
  ram[2440]  = 72;
  ram[2441]  = 72;
  ram[2442]  = 72;
  ram[2443]  = 73;
  ram[2444]  = 73;
  ram[2445]  = 72;
  ram[2446]  = 72;
  ram[2447]  = 73;
  ram[2448]  = 72;
  ram[2449]  = 72;
  ram[2450]  = 72;
  ram[2451]  = 72;
  ram[2452]  = 70;
  ram[2453]  = 70;
  ram[2454]  = 72;
  ram[2455]  = 72;
  ram[2456]  = 73;
  ram[2457]  = 73;
  ram[2458]  = 75;
  ram[2459]  = 73;
  ram[2460]  = 73;
  ram[2461]  = 71;
  ram[2462]  = 72;
  ram[2463]  = 72;
  ram[2464]  = 74;
  ram[2465]  = 73;
  ram[2466]  = 73;
  ram[2467]  = 72;
  ram[2468]  = 70;
  ram[2469]  = 69;
  ram[2470]  = 72;
  ram[2471]  = 74;
  ram[2472]  = 75;
  ram[2473]  = 76;
  ram[2474]  = 77;
  ram[2475]  = 75;
  ram[2476]  = 68;
  ram[2477]  = 68;
  ram[2478]  = 75;
  ram[2479]  = 77;
  ram[2480]  = 72;
  ram[2481]  = 71;
  ram[2482]  = 73;
  ram[2483]  = 73;
  ram[2484]  = 73;
  ram[2485]  = 72;
  ram[2486]  = 70;
  ram[2487]  = 70;
  ram[2488]  = 70;
  ram[2489]  = 70;
  ram[2490]  = 70;
  ram[2491]  = 70;
  ram[2492]  = 70;
  ram[2493]  = 69;
  ram[2494]  = 68;
  ram[2495]  = 68;
  ram[2496]  = 68;
  ram[2497]  = 68;
  ram[2498]  = 69;
  ram[2499]  = 69;
  ram[2500]  = 69;
  ram[2501]  = 68;
  ram[2502]  = 69;
  ram[2503]  = 68;
  ram[2504]  = 70;
  ram[2505]  = 69;
  ram[2506]  = 69;
  ram[2507]  = 70;
  ram[2508]  = 70;
  ram[2509]  = 70;
  ram[2510]  = 72;
  ram[2511]  = 71;
  ram[2512]  = 69;
  ram[2513]  = 69;
  ram[2514]  = 67;
  ram[2515]  = 65;
  ram[2516]  = 63;
  ram[2517]  = 61;
  ram[2518]  = 61;
  ram[2519]  = 62;
  ram[2520]  = 63;
  ram[2521]  = 63;
  ram[2522]  = 66;
  ram[2523]  = 66;
  ram[2524]  = 66;
  ram[2525]  = 64;
  ram[2526]  = 65;
  ram[2527]  = 65;
  ram[2528]  = 66;
  ram[2529]  = 65;
  ram[2530]  = 64;
  ram[2531]  = 63;
  ram[2532]  = 62;
  ram[2533]  = 61;
  ram[2534]  = 65;
  ram[2535]  = 67;
  ram[2536]  = 67;
  ram[2537]  = 68;
  ram[2538]  = 70;
  ram[2539]  = 67;
  ram[2540]  = 60;
  ram[2541]  = 60;
  ram[2542]  = 69;
  ram[2543]  = 73;
  ram[2544]  = 68;
  ram[2545]  = 67;
  ram[2546]  = 68;
  ram[2547]  = 69;
  ram[2548]  = 70;
  ram[2549]  = 70;
  ram[2550]  = 70;
  ram[2551]  = 68;
  ram[2552]  = 68;
  ram[2553]  = 67;
  ram[2554]  = 67;
  ram[2555]  = 67;
  ram[2556]  = 67;
  ram[2557]  = 66;
  ram[2558]  = 65;
  ram[2559]  = 65;
  ram[2560]  = 69;
  ram[2561]  = 69;
  ram[2562]  = 69;
  ram[2563]  = 68;
  ram[2564]  = 68;
  ram[2565]  = 68;
  ram[2566]  = 70;
  ram[2567]  = 70;
  ram[2568]  = 69;
  ram[2569]  = 70;
  ram[2570]  = 70;
  ram[2571]  = 69;
  ram[2572]  = 69;
  ram[2573]  = 69;
  ram[2574]  = 72;
  ram[2575]  = 69;
  ram[2576]  = 63;
  ram[2577]  = 44;
  ram[2578]  = 44;
  ram[2579]  = 37;
  ram[2580]  = 34;
  ram[2581]  = 31;
  ram[2582]  = 32;
  ram[2583]  = 29;
  ram[2584]  = 28;
  ram[2585]  = 30;
  ram[2586]  = 33;
  ram[2587]  = 31;
  ram[2588]  = 34;
  ram[2589]  = 33;
  ram[2590]  = 34;
  ram[2591]  = 35;
  ram[2592]  = 32;
  ram[2593]  = 28;
  ram[2594]  = 34;
  ram[2595]  = 30;
  ram[2596]  = 33;
  ram[2597]  = 32;
  ram[2598]  = 28;
  ram[2599]  = 33;
  ram[2600]  = 26;
  ram[2601]  = 27;
  ram[2602]  = 35;
  ram[2603]  = 30;
  ram[2604]  = 28;
  ram[2605]  = 35;
  ram[2606]  = 39;
  ram[2607]  = 66;
  ram[2608]  = 66;
  ram[2609]  = 69;
  ram[2610]  = 69;
  ram[2611]  = 68;
  ram[2612]  = 69;
  ram[2613]  = 69;
  ram[2614]  = 70;
  ram[2615]  = 67;
  ram[2616]  = 69;
  ram[2617]  = 68;
  ram[2618]  = 68;
  ram[2619]  = 68;
  ram[2620]  = 68;
  ram[2621]  = 67;
  ram[2622]  = 66;
  ram[2623]  = 65;
  ram[2624]  = 70;
  ram[2625]  = 70;
  ram[2626]  = 70;
  ram[2627]  = 70;
  ram[2628]  = 69;
  ram[2629]  = 69;
  ram[2630]  = 69;
  ram[2631]  = 69;
  ram[2632]  = 69;
  ram[2633]  = 69;
  ram[2634]  = 71;
  ram[2635]  = 71;
  ram[2636]  = 71;
  ram[2637]  = 71;
  ram[2638]  = 72;
  ram[2639]  = 67;
  ram[2640]  = 58;
  ram[2641]  = 137;
  ram[2642]  = 131;
  ram[2643]  = 127;
  ram[2644]  = 124;
  ram[2645]  = 115;
  ram[2646]  = 109;
  ram[2647]  = 115;
  ram[2648]  = 113;
  ram[2649]  = 116;
  ram[2650]  = 109;
  ram[2651]  = 118;
  ram[2652]  = 114;
  ram[2653]  = 124;
  ram[2654]  = 117;
  ram[2655]  = 118;
  ram[2656]  = 115;
  ram[2657]  = 118;
  ram[2658]  = 118;
  ram[2659]  = 113;
  ram[2660]  = 119;
  ram[2661]  = 109;
  ram[2662]  = 125;
  ram[2663]  = 108;
  ram[2664]  = 111;
  ram[2665]  = 108;
  ram[2666]  = 113;
  ram[2667]  = 112;
  ram[2668]  = 107;
  ram[2669]  = 102;
  ram[2670]  = 136;
  ram[2671]  = 56;
  ram[2672]  = 64;
  ram[2673]  = 70;
  ram[2674]  = 72;
  ram[2675]  = 68;
  ram[2676]  = 69;
  ram[2677]  = 68;
  ram[2678]  = 69;
  ram[2679]  = 67;
  ram[2680]  = 70;
  ram[2681]  = 68;
  ram[2682]  = 68;
  ram[2683]  = 66;
  ram[2684]  = 68;
  ram[2685]  = 66;
  ram[2686]  = 67;
  ram[2687]  = 65;
  ram[2688]  = 70;
  ram[2689]  = 70;
  ram[2690]  = 70;
  ram[2691]  = 69;
  ram[2692]  = 69;
  ram[2693]  = 69;
  ram[2694]  = 69;
  ram[2695]  = 69;
  ram[2696]  = 69;
  ram[2697]  = 69;
  ram[2698]  = 69;
  ram[2699]  = 70;
  ram[2700]  = 70;
  ram[2701]  = 70;
  ram[2702]  = 72;
  ram[2703]  = 62;
  ram[2704]  = 52;
  ram[2705]  = 195;
  ram[2706]  = 196;
  ram[2707]  = 186;
  ram[2708]  = 178;
  ram[2709]  = 180;
  ram[2710]  = 176;
  ram[2711]  = 172;
  ram[2712]  = 173;
  ram[2713]  = 174;
  ram[2714]  = 170;
  ram[2715]  = 177;
  ram[2716]  = 176;
  ram[2717]  = 181;
  ram[2718]  = 177;
  ram[2719]  = 177;
  ram[2720]  = 178;
  ram[2721]  = 174;
  ram[2722]  = 177;
  ram[2723]  = 175;
  ram[2724]  = 175;
  ram[2725]  = 177;
  ram[2726]  = 179;
  ram[2727]  = 182;
  ram[2728]  = 171;
  ram[2729]  = 166;
  ram[2730]  = 177;
  ram[2731]  = 175;
  ram[2732]  = 158;
  ram[2733]  = 149;
  ram[2734]  = 158;
  ram[2735]  = 44;
  ram[2736]  = 58;
  ram[2737]  = 68;
  ram[2738]  = 70;
  ram[2739]  = 69;
  ram[2740]  = 69;
  ram[2741]  = 68;
  ram[2742]  = 69;
  ram[2743]  = 69;
  ram[2744]  = 70;
  ram[2745]  = 69;
  ram[2746]  = 68;
  ram[2747]  = 66;
  ram[2748]  = 68;
  ram[2749]  = 66;
  ram[2750]  = 69;
  ram[2751]  = 67;
  ram[2752]  = 70;
  ram[2753]  = 68;
  ram[2754]  = 70;
  ram[2755]  = 68;
  ram[2756]  = 68;
  ram[2757]  = 66;
  ram[2758]  = 67;
  ram[2759]  = 67;
  ram[2760]  = 67;
  ram[2761]  = 67;
  ram[2762]  = 67;
  ram[2763]  = 69;
  ram[2764]  = 70;
  ram[2765]  = 70;
  ram[2766]  = 72;
  ram[2767]  = 62;
  ram[2768]  = 46;
  ram[2769]  = 71;
  ram[2770]  = 54;
  ram[2771]  = 55;
  ram[2772]  = 54;
  ram[2773]  = 44;
  ram[2774]  = 44;
  ram[2775]  = 45;
  ram[2776]  = 41;
  ram[2777]  = 45;
  ram[2778]  = 38;
  ram[2779]  = 53;
  ram[2780]  = 40;
  ram[2781]  = 52;
  ram[2782]  = 41;
  ram[2783]  = 46;
  ram[2784]  = 45;
  ram[2785]  = 51;
  ram[2786]  = 44;
  ram[2787]  = 37;
  ram[2788]  = 48;
  ram[2789]  = 41;
  ram[2790]  = 54;
  ram[2791]  = 45;
  ram[2792]  = 51;
  ram[2793]  = 39;
  ram[2794]  = 53;
  ram[2795]  = 32;
  ram[2796]  = 20;
  ram[2797]  = 122;
  ram[2798]  = 147;
  ram[2799]  = 29;
  ram[2800]  = 51;
  ram[2801]  = 66;
  ram[2802]  = 68;
  ram[2803]  = 67;
  ram[2804]  = 66;
  ram[2805]  = 67;
  ram[2806]  = 68;
  ram[2807]  = 69;
  ram[2808]  = 68;
  ram[2809]  = 68;
  ram[2810]  = 67;
  ram[2811]  = 67;
  ram[2812]  = 67;
  ram[2813]  = 67;
  ram[2814]  = 67;
  ram[2815]  = 68;
  ram[2816]  = 72;
  ram[2817]  = 70;
  ram[2818]  = 72;
  ram[2819]  = 69;
  ram[2820]  = 69;
  ram[2821]  = 67;
  ram[2822]  = 69;
  ram[2823]  = 69;
  ram[2824]  = 68;
  ram[2825]  = 69;
  ram[2826]  = 69;
  ram[2827]  = 71;
  ram[2828]  = 71;
  ram[2829]  = 70;
  ram[2830]  = 72;
  ram[2831]  = 69;
  ram[2832]  = 66;
  ram[2833]  = 49;
  ram[2834]  = 53;
  ram[2835]  = 48;
  ram[2836]  = 45;
  ram[2837]  = 38;
  ram[2838]  = 43;
  ram[2839]  = 40;
  ram[2840]  = 43;
  ram[2841]  = 41;
  ram[2842]  = 45;
  ram[2843]  = 43;
  ram[2844]  = 43;
  ram[2845]  = 40;
  ram[2846]  = 44;
  ram[2847]  = 40;
  ram[2848]  = 51;
  ram[2849]  = 42;
  ram[2850]  = 42;
  ram[2851]  = 40;
  ram[2852]  = 38;
  ram[2853]  = 43;
  ram[2854]  = 51;
  ram[2855]  = 48;
  ram[2856]  = 47;
  ram[2857]  = 48;
  ram[2858]  = 47;
  ram[2859]  = 33;
  ram[2860]  = 0;
  ram[2861]  = 140;
  ram[2862]  = 150;
  ram[2863]  = 30;
  ram[2864]  = 53;
  ram[2865]  = 68;
  ram[2866]  = 70;
  ram[2867]  = 69;
  ram[2868]  = 68;
  ram[2869]  = 68;
  ram[2870]  = 69;
  ram[2871]  = 69;
  ram[2872]  = 68;
  ram[2873]  = 68;
  ram[2874]  = 69;
  ram[2875]  = 69;
  ram[2876]  = 69;
  ram[2877]  = 68;
  ram[2878]  = 67;
  ram[2879]  = 67;
  ram[2880]  = 73;
  ram[2881]  = 73;
  ram[2882]  = 72;
  ram[2883]  = 72;
  ram[2884]  = 72;
  ram[2885]  = 69;
  ram[2886]  = 69;
  ram[2887]  = 69;
  ram[2888]  = 70;
  ram[2889]  = 71;
  ram[2890]  = 73;
  ram[2891]  = 72;
  ram[2892]  = 73;
  ram[2893]  = 72;
  ram[2894]  = 72;
  ram[2895]  = 72;
  ram[2896]  = 74;
  ram[2897]  = 69;
  ram[2898]  = 73;
  ram[2899]  = 69;
  ram[2900]  = 70;
  ram[2901]  = 68;
  ram[2902]  = 71;
  ram[2903]  = 70;
  ram[2904]  = 72;
  ram[2905]  = 72;
  ram[2906]  = 72;
  ram[2907]  = 73;
  ram[2908]  = 65;
  ram[2909]  = 72;
  ram[2910]  = 70;
  ram[2911]  = 68;
  ram[2912]  = 66;
  ram[2913]  = 70;
  ram[2914]  = 66;
  ram[2915]  = 66;
  ram[2916]  = 65;
  ram[2917]  = 62;
  ram[2918]  = 69;
  ram[2919]  = 70;
  ram[2920]  = 65;
  ram[2921]  = 60;
  ram[2922]  = 61;
  ram[2923]  = 36;
  ram[2924]  = 6;
  ram[2925]  = 135;
  ram[2926]  = 150;
  ram[2927]  = 30;
  ram[2928]  = 53;
  ram[2929]  = 68;
  ram[2930]  = 70;
  ram[2931]  = 69;
  ram[2932]  = 69;
  ram[2933]  = 69;
  ram[2934]  = 70;
  ram[2935]  = 70;
  ram[2936]  = 69;
  ram[2937]  = 69;
  ram[2938]  = 72;
  ram[2939]  = 72;
  ram[2940]  = 72;
  ram[2941]  = 71;
  ram[2942]  = 70;
  ram[2943]  = 70;
  ram[2944]  = 74;
  ram[2945]  = 74;
  ram[2946]  = 74;
  ram[2947]  = 71;
  ram[2948]  = 71;
  ram[2949]  = 71;
  ram[2950]  = 70;
  ram[2951]  = 70;
  ram[2952]  = 72;
  ram[2953]  = 71;
  ram[2954]  = 73;
  ram[2955]  = 72;
  ram[2956]  = 74;
  ram[2957]  = 73;
  ram[2958]  = 73;
  ram[2959]  = 71;
  ram[2960]  = 66;
  ram[2961]  = 74;
  ram[2962]  = 70;
  ram[2963]  = 68;
  ram[2964]  = 72;
  ram[2965]  = 73;
  ram[2966]  = 71;
  ram[2967]  = 71;
  ram[2968]  = 75;
  ram[2969]  = 71;
  ram[2970]  = 76;
  ram[2971]  = 70;
  ram[2972]  = 73;
  ram[2973]  = 69;
  ram[2974]  = 69;
  ram[2975]  = 57;
  ram[2976]  = 84;
  ram[2977]  = 81;
  ram[2978]  = 65;
  ram[2979]  = 70;
  ram[2980]  = 67;
  ram[2981]  = 67;
  ram[2982]  = 61;
  ram[2983]  = 57;
  ram[2984]  = 50;
  ram[2985]  = 38;
  ram[2986]  = 37;
  ram[2987]  = 30;
  ram[2988]  = 0;
  ram[2989]  = 131;
  ram[2990]  = 156;
  ram[2991]  = 26;
  ram[2992]  = 54;
  ram[2993]  = 68;
  ram[2994]  = 70;
  ram[2995]  = 70;
  ram[2996]  = 71;
  ram[2997]  = 71;
  ram[2998]  = 72;
  ram[2999]  = 71;
  ram[3000]  = 71;
  ram[3001]  = 71;
  ram[3002]  = 73;
  ram[3003]  = 73;
  ram[3004]  = 73;
  ram[3005]  = 73;
  ram[3006]  = 72;
  ram[3007]  = 72;
  ram[3008]  = 75;
  ram[3009]  = 72;
  ram[3010]  = 74;
  ram[3011]  = 72;
  ram[3012]  = 71;
  ram[3013]  = 71;
  ram[3014]  = 71;
  ram[3015]  = 71;
  ram[3016]  = 71;
  ram[3017]  = 70;
  ram[3018]  = 70;
  ram[3019]  = 72;
  ram[3020]  = 72;
  ram[3021]  = 73;
  ram[3022]  = 73;
  ram[3023]  = 70;
  ram[3024]  = 69;
  ram[3025]  = 65;
  ram[3026]  = 66;
  ram[3027]  = 70;
  ram[3028]  = 69;
  ram[3029]  = 71;
  ram[3030]  = 73;
  ram[3031]  = 75;
  ram[3032]  = 76;
  ram[3033]  = 73;
  ram[3034]  = 74;
  ram[3035]  = 73;
  ram[3036]  = 70;
  ram[3037]  = 71;
  ram[3038]  = 61;
  ram[3039]  = 41;
  ram[3040]  = 255;
  ram[3041]  = 255;
  ram[3042]  = 43;
  ram[3043]  = 74;
  ram[3044]  = 76;
  ram[3045]  = 67;
  ram[3046]  = 51;
  ram[3047]  = 137;
  ram[3048]  = 194;
  ram[3049]  = 161;
  ram[3050]  = 167;
  ram[3051]  = 157;
  ram[3052]  = 145;
  ram[3053]  = 135;
  ram[3054]  = 160;
  ram[3055]  = 40;
  ram[3056]  = 58;
  ram[3057]  = 70;
  ram[3058]  = 71;
  ram[3059]  = 69;
  ram[3060]  = 71;
  ram[3061]  = 69;
  ram[3062]  = 70;
  ram[3063]  = 69;
  ram[3064]  = 70;
  ram[3065]  = 70;
  ram[3066]  = 70;
  ram[3067]  = 70;
  ram[3068]  = 70;
  ram[3069]  = 70;
  ram[3070]  = 71;
  ram[3071]  = 71;
  ram[3072]  = 74;
  ram[3073]  = 73;
  ram[3074]  = 75;
  ram[3075]  = 74;
  ram[3076]  = 74;
  ram[3077]  = 74;
  ram[3078]  = 73;
  ram[3079]  = 73;
  ram[3080]  = 74;
  ram[3081]  = 74;
  ram[3082]  = 74;
  ram[3083]  = 75;
  ram[3084]  = 75;
  ram[3085]  = 75;
  ram[3086]  = 75;
  ram[3087]  = 74;
  ram[3088]  = 71;
  ram[3089]  = 70;
  ram[3090]  = 69;
  ram[3091]  = 70;
  ram[3092]  = 71;
  ram[3093]  = 74;
  ram[3094]  = 73;
  ram[3095]  = 71;
  ram[3096]  = 74;
  ram[3097]  = 73;
  ram[3098]  = 73;
  ram[3099]  = 74;
  ram[3100]  = 71;
  ram[3101]  = 74;
  ram[3102]  = 71;
  ram[3103]  = 43;
  ram[3104]  = 233;
  ram[3105]  = 219;
  ram[3106]  = 42;
  ram[3107]  = 76;
  ram[3108]  = 80;
  ram[3109]  = 79;
  ram[3110]  = 55;
  ram[3111]  = 120;
  ram[3112]  = 174;
  ram[3113]  = 154;
  ram[3114]  = 146;
  ram[3115]  = 137;
  ram[3116]  = 140;
  ram[3117]  = 145;
  ram[3118]  = 148;
  ram[3119]  = 50;
  ram[3120]  = 63;
  ram[3121]  = 71;
  ram[3122]  = 71;
  ram[3123]  = 70;
  ram[3124]  = 72;
  ram[3125]  = 71;
  ram[3126]  = 74;
  ram[3127]  = 74;
  ram[3128]  = 74;
  ram[3129]  = 74;
  ram[3130]  = 74;
  ram[3131]  = 73;
  ram[3132]  = 73;
  ram[3133]  = 73;
  ram[3134]  = 73;
  ram[3135]  = 72;
  ram[3136]  = 75;
  ram[3137]  = 75;
  ram[3138]  = 75;
  ram[3139]  = 76;
  ram[3140]  = 76;
  ram[3141]  = 75;
  ram[3142]  = 75;
  ram[3143]  = 75;
  ram[3144]  = 74;
  ram[3145]  = 74;
  ram[3146]  = 74;
  ram[3147]  = 74;
  ram[3148]  = 74;
  ram[3149]  = 74;
  ram[3150]  = 75;
  ram[3151]  = 75;
  ram[3152]  = 73;
  ram[3153]  = 72;
  ram[3154]  = 72;
  ram[3155]  = 72;
  ram[3156]  = 74;
  ram[3157]  = 74;
  ram[3158]  = 73;
  ram[3159]  = 72;
  ram[3160]  = 72;
  ram[3161]  = 72;
  ram[3162]  = 73;
  ram[3163]  = 75;
  ram[3164]  = 71;
  ram[3165]  = 73;
  ram[3166]  = 76;
  ram[3167]  = 61;
  ram[3168]  = 60;
  ram[3169]  = 55;
  ram[3170]  = 71;
  ram[3171]  = 78;
  ram[3172]  = 80;
  ram[3173]  = 82;
  ram[3174]  = 71;
  ram[3175]  = 56;
  ram[3176]  = 32;
  ram[3177]  = 24;
  ram[3178]  = 23;
  ram[3179]  = 16;
  ram[3180]  = 27;
  ram[3181]  = 27;
  ram[3182]  = 43;
  ram[3183]  = 54;
  ram[3184]  = 68;
  ram[3185]  = 73;
  ram[3186]  = 73;
  ram[3187]  = 73;
  ram[3188]  = 73;
  ram[3189]  = 74;
  ram[3190]  = 74;
  ram[3191]  = 74;
  ram[3192]  = 73;
  ram[3193]  = 74;
  ram[3194]  = 74;
  ram[3195]  = 73;
  ram[3196]  = 73;
  ram[3197]  = 73;
  ram[3198]  = 74;
  ram[3199]  = 73;
  ram[3200]  = 75;
  ram[3201]  = 75;
  ram[3202]  = 75;
  ram[3203]  = 75;
  ram[3204]  = 75;
  ram[3205]  = 74;
  ram[3206]  = 74;
  ram[3207]  = 74;
  ram[3208]  = 74;
  ram[3209]  = 73;
  ram[3210]  = 73;
  ram[3211]  = 73;
  ram[3212]  = 74;
  ram[3213]  = 74;
  ram[3214]  = 74;
  ram[3215]  = 74;
  ram[3216]  = 73;
  ram[3217]  = 72;
  ram[3218]  = 72;
  ram[3219]  = 72;
  ram[3220]  = 73;
  ram[3221]  = 74;
  ram[3222]  = 73;
  ram[3223]  = 72;
  ram[3224]  = 71;
  ram[3225]  = 71;
  ram[3226]  = 72;
  ram[3227]  = 74;
  ram[3228]  = 72;
  ram[3229]  = 71;
  ram[3230]  = 76;
  ram[3231]  = 74;
  ram[3232]  = 61;
  ram[3233]  = 68;
  ram[3234]  = 70;
  ram[3235]  = 73;
  ram[3236]  = 76;
  ram[3237]  = 71;
  ram[3238]  = 69;
  ram[3239]  = 63;
  ram[3240]  = 68;
  ram[3241]  = 58;
  ram[3242]  = 61;
  ram[3243]  = 56;
  ram[3244]  = 57;
  ram[3245]  = 67;
  ram[3246]  = 69;
  ram[3247]  = 74;
  ram[3248]  = 73;
  ram[3249]  = 73;
  ram[3250]  = 73;
  ram[3251]  = 73;
  ram[3252]  = 73;
  ram[3253]  = 73;
  ram[3254]  = 74;
  ram[3255]  = 74;
  ram[3256]  = 73;
  ram[3257]  = 74;
  ram[3258]  = 74;
  ram[3259]  = 73;
  ram[3260]  = 74;
  ram[3261]  = 74;
  ram[3262]  = 74;
  ram[3263]  = 73;
  ram[3264]  = 75;
  ram[3265]  = 75;
  ram[3266]  = 75;
  ram[3267]  = 75;
  ram[3268]  = 74;
  ram[3269]  = 74;
  ram[3270]  = 74;
  ram[3271]  = 74;
  ram[3272]  = 74;
  ram[3273]  = 74;
  ram[3274]  = 74;
  ram[3275]  = 74;
  ram[3276]  = 75;
  ram[3277]  = 75;
  ram[3278]  = 75;
  ram[3279]  = 75;
  ram[3280]  = 74;
  ram[3281]  = 73;
  ram[3282]  = 73;
  ram[3283]  = 73;
  ram[3284]  = 74;
  ram[3285]  = 74;
  ram[3286]  = 73;
  ram[3287]  = 72;
  ram[3288]  = 73;
  ram[3289]  = 73;
  ram[3290]  = 71;
  ram[3291]  = 73;
  ram[3292]  = 74;
  ram[3293]  = 73;
  ram[3294]  = 73;
  ram[3295]  = 74;
  ram[3296]  = 78;
  ram[3297]  = 74;
  ram[3298]  = 71;
  ram[3299]  = 76;
  ram[3300]  = 67;
  ram[3301]  = 69;
  ram[3302]  = 75;
  ram[3303]  = 72;
  ram[3304]  = 69;
  ram[3305]  = 76;
  ram[3306]  = 80;
  ram[3307]  = 82;
  ram[3308]  = 78;
  ram[3309]  = 80;
  ram[3310]  = 78;
  ram[3311]  = 78;
  ram[3312]  = 75;
  ram[3313]  = 73;
  ram[3314]  = 73;
  ram[3315]  = 74;
  ram[3316]  = 73;
  ram[3317]  = 74;
  ram[3318]  = 74;
  ram[3319]  = 75;
  ram[3320]  = 74;
  ram[3321]  = 75;
  ram[3322]  = 74;
  ram[3323]  = 74;
  ram[3324]  = 74;
  ram[3325]  = 74;
  ram[3326]  = 74;
  ram[3327]  = 73;
  ram[3328]  = 76;
  ram[3329]  = 76;
  ram[3330]  = 76;
  ram[3331]  = 76;
  ram[3332]  = 76;
  ram[3333]  = 76;
  ram[3334]  = 76;
  ram[3335]  = 76;
  ram[3336]  = 76;
  ram[3337]  = 76;
  ram[3338]  = 76;
  ram[3339]  = 76;
  ram[3340]  = 76;
  ram[3341]  = 76;
  ram[3342]  = 76;
  ram[3343]  = 76;
  ram[3344]  = 76;
  ram[3345]  = 76;
  ram[3346]  = 75;
  ram[3347]  = 76;
  ram[3348]  = 76;
  ram[3349]  = 76;
  ram[3350]  = 76;
  ram[3351]  = 75;
  ram[3352]  = 75;
  ram[3353]  = 77;
  ram[3354]  = 75;
  ram[3355]  = 74;
  ram[3356]  = 76;
  ram[3357]  = 76;
  ram[3358]  = 74;
  ram[3359]  = 76;
  ram[3360]  = 78;
  ram[3361]  = 79;
  ram[3362]  = 79;
  ram[3363]  = 73;
  ram[3364]  = 69;
  ram[3365]  = 72;
  ram[3366]  = 67;
  ram[3367]  = 74;
  ram[3368]  = 77;
  ram[3369]  = 75;
  ram[3370]  = 75;
  ram[3371]  = 82;
  ram[3372]  = 78;
  ram[3373]  = 71;
  ram[3374]  = 77;
  ram[3375]  = 71;
  ram[3376]  = 75;
  ram[3377]  = 75;
  ram[3378]  = 75;
  ram[3379]  = 76;
  ram[3380]  = 76;
  ram[3381]  = 76;
  ram[3382]  = 76;
  ram[3383]  = 77;
  ram[3384]  = 76;
  ram[3385]  = 76;
  ram[3386]  = 76;
  ram[3387]  = 75;
  ram[3388]  = 75;
  ram[3389]  = 75;
  ram[3390]  = 74;
  ram[3391]  = 73;
  ram[3392]  = 76;
  ram[3393]  = 76;
  ram[3394]  = 76;
  ram[3395]  = 76;
  ram[3396]  = 76;
  ram[3397]  = 77;
  ram[3398]  = 77;
  ram[3399]  = 77;
  ram[3400]  = 78;
  ram[3401]  = 78;
  ram[3402]  = 78;
  ram[3403]  = 78;
  ram[3404]  = 78;
  ram[3405]  = 78;
  ram[3406]  = 78;
  ram[3407]  = 77;
  ram[3408]  = 76;
  ram[3409]  = 76;
  ram[3410]  = 75;
  ram[3411]  = 76;
  ram[3412]  = 76;
  ram[3413]  = 76;
  ram[3414]  = 75;
  ram[3415]  = 75;
  ram[3416]  = 73;
  ram[3417]  = 76;
  ram[3418]  = 78;
  ram[3419]  = 74;
  ram[3420]  = 74;
  ram[3421]  = 76;
  ram[3422]  = 75;
  ram[3423]  = 80;
  ram[3424]  = 85;
  ram[3425]  = 80;
  ram[3426]  = 74;
  ram[3427]  = 84;
  ram[3428]  = 71;
  ram[3429]  = 74;
  ram[3430]  = 76;
  ram[3431]  = 72;
  ram[3432]  = 71;
  ram[3433]  = 80;
  ram[3434]  = 79;
  ram[3435]  = 72;
  ram[3436]  = 79;
  ram[3437]  = 71;
  ram[3438]  = 67;
  ram[3439]  = 78;
  ram[3440]  = 77;
  ram[3441]  = 77;
  ram[3442]  = 77;
  ram[3443]  = 76;
  ram[3444]  = 76;
  ram[3445]  = 76;
  ram[3446]  = 76;
  ram[3447]  = 76;
  ram[3448]  = 77;
  ram[3449]  = 78;
  ram[3450]  = 78;
  ram[3451]  = 77;
  ram[3452]  = 76;
  ram[3453]  = 76;
  ram[3454]  = 75;
  ram[3455]  = 74;
  ram[3456]  = 76;
  ram[3457]  = 76;
  ram[3458]  = 76;
  ram[3459]  = 76;
  ram[3460]  = 77;
  ram[3461]  = 77;
  ram[3462]  = 78;
  ram[3463]  = 78;
  ram[3464]  = 79;
  ram[3465]  = 79;
  ram[3466]  = 79;
  ram[3467]  = 79;
  ram[3468]  = 79;
  ram[3469]  = 78;
  ram[3470]  = 78;
  ram[3471]  = 77;
  ram[3472]  = 76;
  ram[3473]  = 76;
  ram[3474]  = 75;
  ram[3475]  = 75;
  ram[3476]  = 76;
  ram[3477]  = 75;
  ram[3478]  = 75;
  ram[3479]  = 74;
  ram[3480]  = 74;
  ram[3481]  = 74;
  ram[3482]  = 78;
  ram[3483]  = 76;
  ram[3484]  = 74;
  ram[3485]  = 77;
  ram[3486]  = 76;
  ram[3487]  = 79;
  ram[3488]  = 77;
  ram[3489]  = 76;
  ram[3490]  = 84;
  ram[3491]  = 80;
  ram[3492]  = 75;
  ram[3493]  = 76;
  ram[3494]  = 81;
  ram[3495]  = 74;
  ram[3496]  = 85;
  ram[3497]  = 70;
  ram[3498]  = 74;
  ram[3499]  = 75;
  ram[3500]  = 72;
  ram[3501]  = 72;
  ram[3502]  = 77;
  ram[3503]  = 76;
  ram[3504]  = 78;
  ram[3505]  = 79;
  ram[3506]  = 79;
  ram[3507]  = 79;
  ram[3508]  = 76;
  ram[3509]  = 76;
  ram[3510]  = 76;
  ram[3511]  = 76;
  ram[3512]  = 78;
  ram[3513]  = 79;
  ram[3514]  = 79;
  ram[3515]  = 78;
  ram[3516]  = 79;
  ram[3517]  = 79;
  ram[3518]  = 78;
  ram[3519]  = 77;
  ram[3520]  = 78;
  ram[3521]  = 77;
  ram[3522]  = 77;
  ram[3523]  = 78;
  ram[3524]  = 78;
  ram[3525]  = 79;
  ram[3526]  = 79;
  ram[3527]  = 80;
  ram[3528]  = 79;
  ram[3529]  = 79;
  ram[3530]  = 79;
  ram[3531]  = 79;
  ram[3532]  = 79;
  ram[3533]  = 78;
  ram[3534]  = 77;
  ram[3535]  = 77;
  ram[3536]  = 78;
  ram[3537]  = 77;
  ram[3538]  = 77;
  ram[3539]  = 77;
  ram[3540]  = 77;
  ram[3541]  = 77;
  ram[3542]  = 76;
  ram[3543]  = 76;
  ram[3544]  = 78;
  ram[3545]  = 74;
  ram[3546]  = 79;
  ram[3547]  = 79;
  ram[3548]  = 79;
  ram[3549]  = 80;
  ram[3550]  = 77;
  ram[3551]  = 77;
  ram[3552]  = 77;
  ram[3553]  = 84;
  ram[3554]  = 75;
  ram[3555]  = 81;
  ram[3556]  = 83;
  ram[3557]  = 79;
  ram[3558]  = 77;
  ram[3559]  = 77;
  ram[3560]  = 75;
  ram[3561]  = 81;
  ram[3562]  = 77;
  ram[3563]  = 75;
  ram[3564]  = 76;
  ram[3565]  = 80;
  ram[3566]  = 82;
  ram[3567]  = 78;
  ram[3568]  = 80;
  ram[3569]  = 80;
  ram[3570]  = 80;
  ram[3571]  = 80;
  ram[3572]  = 78;
  ram[3573]  = 78;
  ram[3574]  = 78;
  ram[3575]  = 79;
  ram[3576]  = 78;
  ram[3577]  = 79;
  ram[3578]  = 80;
  ram[3579]  = 79;
  ram[3580]  = 80;
  ram[3581]  = 80;
  ram[3582]  = 79;
  ram[3583]  = 77;
  ram[3584]  = 79;
  ram[3585]  = 79;
  ram[3586]  = 79;
  ram[3587]  = 78;
  ram[3588]  = 78;
  ram[3589]  = 78;
  ram[3590]  = 78;
  ram[3591]  = 77;
  ram[3592]  = 77;
  ram[3593]  = 77;
  ram[3594]  = 77;
  ram[3595]  = 77;
  ram[3596]  = 77;
  ram[3597]  = 77;
  ram[3598]  = 77;
  ram[3599]  = 77;
  ram[3600]  = 76;
  ram[3601]  = 76;
  ram[3602]  = 76;
  ram[3603]  = 77;
  ram[3604]  = 77;
  ram[3605]  = 77;
  ram[3606]  = 77;
  ram[3607]  = 77;
  ram[3608]  = 77;
  ram[3609]  = 77;
  ram[3610]  = 77;
  ram[3611]  = 77;
  ram[3612]  = 77;
  ram[3613]  = 77;
  ram[3614]  = 77;
  ram[3615]  = 77;
  ram[3616]  = 80;
  ram[3617]  = 80;
  ram[3618]  = 79;
  ram[3619]  = 77;
  ram[3620]  = 79;
  ram[3621]  = 79;
  ram[3622]  = 79;
  ram[3623]  = 79;
  ram[3624]  = 79;
  ram[3625]  = 79;
  ram[3626]  = 81;
  ram[3627]  = 81;
  ram[3628]  = 82;
  ram[3629]  = 84;
  ram[3630]  = 84;
  ram[3631]  = 82;
  ram[3632]  = 83;
  ram[3633]  = 81;
  ram[3634]  = 81;
  ram[3635]  = 81;
  ram[3636]  = 78;
  ram[3637]  = 78;
  ram[3638]  = 78;
  ram[3639]  = 78;
  ram[3640]  = 79;
  ram[3641]  = 79;
  ram[3642]  = 79;
  ram[3643]  = 79;
  ram[3644]  = 80;
  ram[3645]  = 79;
  ram[3646]  = 79;
  ram[3647]  = 78;
  ram[3648]  = 78;
  ram[3649]  = 79;
  ram[3650]  = 79;
  ram[3651]  = 78;
  ram[3652]  = 78;
  ram[3653]  = 79;
  ram[3654]  = 79;
  ram[3655]  = 78;
  ram[3656]  = 80;
  ram[3657]  = 80;
  ram[3658]  = 80;
  ram[3659]  = 80;
  ram[3660]  = 80;
  ram[3661]  = 80;
  ram[3662]  = 80;
  ram[3663]  = 80;
  ram[3664]  = 80;
  ram[3665]  = 80;
  ram[3666]  = 80;
  ram[3667]  = 80;
  ram[3668]  = 80;
  ram[3669]  = 80;
  ram[3670]  = 80;
  ram[3671]  = 80;
  ram[3672]  = 79;
  ram[3673]  = 79;
  ram[3674]  = 79;
  ram[3675]  = 79;
  ram[3676]  = 79;
  ram[3677]  = 79;
  ram[3678]  = 79;
  ram[3679]  = 79;
  ram[3680]  = 81;
  ram[3681]  = 81;
  ram[3682]  = 79;
  ram[3683]  = 79;
  ram[3684]  = 79;
  ram[3685]  = 79;
  ram[3686]  = 78;
  ram[3687]  = 80;
  ram[3688]  = 81;
  ram[3689]  = 83;
  ram[3690]  = 85;
  ram[3691]  = 85;
  ram[3692]  = 85;
  ram[3693]  = 85;
  ram[3694]  = 86;
  ram[3695]  = 84;
  ram[3696]  = 82;
  ram[3697]  = 82;
  ram[3698]  = 82;
  ram[3699]  = 82;
  ram[3700]  = 80;
  ram[3701]  = 80;
  ram[3702]  = 80;
  ram[3703]  = 80;
  ram[3704]  = 79;
  ram[3705]  = 79;
  ram[3706]  = 79;
  ram[3707]  = 79;
  ram[3708]  = 80;
  ram[3709]  = 79;
  ram[3710]  = 79;
  ram[3711]  = 78;
  ram[3712]  = 79;
  ram[3713]  = 79;
  ram[3714]  = 79;
  ram[3715]  = 78;
  ram[3716]  = 79;
  ram[3717]  = 80;
  ram[3718]  = 80;
  ram[3719]  = 80;
  ram[3720]  = 80;
  ram[3721]  = 80;
  ram[3722]  = 80;
  ram[3723]  = 80;
  ram[3724]  = 79;
  ram[3725]  = 79;
  ram[3726]  = 79;
  ram[3727]  = 79;
  ram[3728]  = 79;
  ram[3729]  = 79;
  ram[3730]  = 79;
  ram[3731]  = 79;
  ram[3732]  = 79;
  ram[3733]  = 79;
  ram[3734]  = 79;
  ram[3735]  = 79;
  ram[3736]  = 79;
  ram[3737]  = 79;
  ram[3738]  = 79;
  ram[3739]  = 79;
  ram[3740]  = 79;
  ram[3741]  = 79;
  ram[3742]  = 79;
  ram[3743]  = 79;
  ram[3744]  = 81;
  ram[3745]  = 81;
  ram[3746]  = 79;
  ram[3747]  = 79;
  ram[3748]  = 78;
  ram[3749]  = 77;
  ram[3750]  = 77;
  ram[3751]  = 78;
  ram[3752]  = 79;
  ram[3753]  = 79;
  ram[3754]  = 81;
  ram[3755]  = 81;
  ram[3756]  = 79;
  ram[3757]  = 79;
  ram[3758]  = 79;
  ram[3759]  = 80;
  ram[3760]  = 81;
  ram[3761]  = 81;
  ram[3762]  = 81;
  ram[3763]  = 81;
  ram[3764]  = 79;
  ram[3765]  = 79;
  ram[3766]  = 79;
  ram[3767]  = 79;
  ram[3768]  = 79;
  ram[3769]  = 79;
  ram[3770]  = 79;
  ram[3771]  = 79;
  ram[3772]  = 80;
  ram[3773]  = 79;
  ram[3774]  = 79;
  ram[3775]  = 78;
  ram[3776]  = 80;
  ram[3777]  = 80;
  ram[3778]  = 80;
  ram[3779]  = 79;
  ram[3780]  = 79;
  ram[3781]  = 80;
  ram[3782]  = 80;
  ram[3783]  = 80;
  ram[3784]  = 81;
  ram[3785]  = 80;
  ram[3786]  = 80;
  ram[3787]  = 80;
  ram[3788]  = 80;
  ram[3789]  = 80;
  ram[3790]  = 80;
  ram[3791]  = 80;
  ram[3792]  = 80;
  ram[3793]  = 80;
  ram[3794]  = 80;
  ram[3795]  = 80;
  ram[3796]  = 80;
  ram[3797]  = 80;
  ram[3798]  = 80;
  ram[3799]  = 80;
  ram[3800]  = 81;
  ram[3801]  = 81;
  ram[3802]  = 81;
  ram[3803]  = 81;
  ram[3804]  = 81;
  ram[3805]  = 80;
  ram[3806]  = 80;
  ram[3807]  = 80;
  ram[3808]  = 81;
  ram[3809]  = 81;
  ram[3810]  = 81;
  ram[3811]  = 80;
  ram[3812]  = 79;
  ram[3813]  = 79;
  ram[3814]  = 79;
  ram[3815]  = 79;
  ram[3816]  = 80;
  ram[3817]  = 80;
  ram[3818]  = 80;
  ram[3819]  = 80;
  ram[3820]  = 81;
  ram[3821]  = 80;
  ram[3822]  = 81;
  ram[3823]  = 81;
  ram[3824]  = 83;
  ram[3825]  = 83;
  ram[3826]  = 82;
  ram[3827]  = 82;
  ram[3828]  = 80;
  ram[3829]  = 80;
  ram[3830]  = 80;
  ram[3831]  = 80;
  ram[3832]  = 79;
  ram[3833]  = 79;
  ram[3834]  = 79;
  ram[3835]  = 79;
  ram[3836]  = 80;
  ram[3837]  = 79;
  ram[3838]  = 79;
  ram[3839]  = 78;
  ram[3840]  = 81;
  ram[3841]  = 81;
  ram[3842]  = 80;
  ram[3843]  = 79;
  ram[3844]  = 79;
  ram[3845]  = 79;
  ram[3846]  = 79;
  ram[3847]  = 79;
  ram[3848]  = 79;
  ram[3849]  = 79;
  ram[3850]  = 79;
  ram[3851]  = 79;
  ram[3852]  = 79;
  ram[3853]  = 79;
  ram[3854]  = 79;
  ram[3855]  = 79;
  ram[3856]  = 79;
  ram[3857]  = 79;
  ram[3858]  = 79;
  ram[3859]  = 79;
  ram[3860]  = 79;
  ram[3861]  = 79;
  ram[3862]  = 80;
  ram[3863]  = 80;
  ram[3864]  = 79;
  ram[3865]  = 79;
  ram[3866]  = 79;
  ram[3867]  = 79;
  ram[3868]  = 79;
  ram[3869]  = 79;
  ram[3870]  = 79;
  ram[3871]  = 78;
  ram[3872]  = 78;
  ram[3873]  = 76;
  ram[3874]  = 79;
  ram[3875]  = 79;
  ram[3876]  = 81;
  ram[3877]  = 81;
  ram[3878]  = 81;
  ram[3879]  = 79;
  ram[3880]  = 79;
  ram[3881]  = 79;
  ram[3882]  = 79;
  ram[3883]  = 79;
  ram[3884]  = 79;
  ram[3885]  = 81;
  ram[3886]  = 83;
  ram[3887]  = 83;
  ram[3888]  = 81;
  ram[3889]  = 81;
  ram[3890]  = 79;
  ram[3891]  = 78;
  ram[3892]  = 78;
  ram[3893]  = 78;
  ram[3894]  = 78;
  ram[3895]  = 79;
  ram[3896]  = 79;
  ram[3897]  = 79;
  ram[3898]  = 79;
  ram[3899]  = 79;
  ram[3900]  = 78;
  ram[3901]  = 78;
  ram[3902]  = 79;
  ram[3903]  = 78;
  ram[3904]  = 80;
  ram[3905]  = 81;
  ram[3906]  = 80;
  ram[3907]  = 79;
  ram[3908]  = 78;
  ram[3909]  = 79;
  ram[3910]  = 79;
  ram[3911]  = 78;
  ram[3912]  = 78;
  ram[3913]  = 78;
  ram[3914]  = 78;
  ram[3915]  = 78;
  ram[3916]  = 78;
  ram[3917]  = 78;
  ram[3918]  = 78;
  ram[3919]  = 78;
  ram[3920]  = 77;
  ram[3921]  = 77;
  ram[3922]  = 77;
  ram[3923]  = 78;
  ram[3924]  = 78;
  ram[3925]  = 78;
  ram[3926]  = 78;
  ram[3927]  = 78;
  ram[3928]  = 78;
  ram[3929]  = 77;
  ram[3930]  = 77;
  ram[3931]  = 77;
  ram[3932]  = 77;
  ram[3933]  = 77;
  ram[3934]  = 77;
  ram[3935]  = 76;
  ram[3936]  = 74;
  ram[3937]  = 74;
  ram[3938]  = 76;
  ram[3939]  = 77;
  ram[3940]  = 79;
  ram[3941]  = 79;
  ram[3942]  = 79;
  ram[3943]  = 77;
  ram[3944]  = 77;
  ram[3945]  = 77;
  ram[3946]  = 77;
  ram[3947]  = 77;
  ram[3948]  = 77;
  ram[3949]  = 79;
  ram[3950]  = 81;
  ram[3951]  = 81;
  ram[3952]  = 79;
  ram[3953]  = 79;
  ram[3954]  = 77;
  ram[3955]  = 77;
  ram[3956]  = 77;
  ram[3957]  = 77;
  ram[3958]  = 77;
  ram[3959]  = 77;
  ram[3960]  = 79;
  ram[3961]  = 79;
  ram[3962]  = 79;
  ram[3963]  = 79;
  ram[3964]  = 78;
  ram[3965]  = 78;
  ram[3966]  = 79;
  ram[3967]  = 78;
  ram[3968]  = 78;
  ram[3969]  = 79;
  ram[3970]  = 79;
  ram[3971]  = 78;
  ram[3972]  = 78;
  ram[3973]  = 79;
  ram[3974]  = 79;
  ram[3975]  = 79;
  ram[3976]  = 81;
  ram[3977]  = 81;
  ram[3978]  = 81;
  ram[3979]  = 81;
  ram[3980]  = 81;
  ram[3981]  = 81;
  ram[3982]  = 81;
  ram[3983]  = 81;
  ram[3984]  = 79;
  ram[3985]  = 79;
  ram[3986]  = 80;
  ram[3987]  = 80;
  ram[3988]  = 80;
  ram[3989]  = 80;
  ram[3990]  = 80;
  ram[3991]  = 80;
  ram[3992]  = 80;
  ram[3993]  = 80;
  ram[3994]  = 80;
  ram[3995]  = 80;
  ram[3996]  = 80;
  ram[3997]  = 80;
  ram[3998]  = 80;
  ram[3999]  = 80;
  ram[4000]  = 79;
  ram[4001]  = 79;
  ram[4002]  = 80;
  ram[4003]  = 80;
  ram[4004]  = 80;
  ram[4005]  = 80;
  ram[4006]  = 80;
  ram[4007]  = 79;
  ram[4008]  = 79;
  ram[4009]  = 79;
  ram[4010]  = 79;
  ram[4011]  = 79;
  ram[4012]  = 78;
  ram[4013]  = 78;
  ram[4014]  = 79;
  ram[4015]  = 79;
  ram[4016]  = 80;
  ram[4017]  = 80;
  ram[4018]  = 80;
  ram[4019]  = 80;
  ram[4020]  = 80;
  ram[4021]  = 80;
  ram[4022]  = 79;
  ram[4023]  = 79;
  ram[4024]  = 78;
  ram[4025]  = 78;
  ram[4026]  = 79;
  ram[4027]  = 79;
  ram[4028]  = 78;
  ram[4029]  = 78;
  ram[4030]  = 77;
  ram[4031]  = 76;
  ram[4032]  = 76;
  ram[4033]  = 77;
  ram[4034]  = 78;
  ram[4035]  = 78;
  ram[4036]  = 79;
  ram[4037]  = 80;
  ram[4038]  = 80;
  ram[4039]  = 79;
  ram[4040]  = 78;
  ram[4041]  = 78;
  ram[4042]  = 78;
  ram[4043]  = 78;
  ram[4044]  = 78;
  ram[4045]  = 78;
  ram[4046]  = 78;
  ram[4047]  = 78;
  ram[4048]  = 78;
  ram[4049]  = 78;
  ram[4050]  = 78;
  ram[4051]  = 78;
  ram[4052]  = 78;
  ram[4053]  = 78;
  ram[4054]  = 78;
  ram[4055]  = 78;
  ram[4056]  = 78;
  ram[4057]  = 78;
  ram[4058]  = 78;
  ram[4059]  = 78;
  ram[4060]  = 78;
  ram[4061]  = 78;
  ram[4062]  = 78;
  ram[4063]  = 78;
  ram[4064]  = 78;
  ram[4065]  = 78;
  ram[4066]  = 78;
  ram[4067]  = 78;
  ram[4068]  = 78;
  ram[4069]  = 78;
  ram[4070]  = 77;
  ram[4071]  = 77;
  ram[4072]  = 77;
  ram[4073]  = 77;
  ram[4074]  = 77;
  ram[4075]  = 77;
  ram[4076]  = 75;
  ram[4077]  = 75;
  ram[4078]  = 73;
  ram[4079]  = 75;
  ram[4080]  = 78;
  ram[4081]  = 79;
  ram[4082]  = 78;
  ram[4083]  = 78;
  ram[4084]  = 78;
  ram[4085]  = 79;
  ram[4086]  = 78;
  ram[4087]  = 78;
  ram[4088]  = 78;
  ram[4089]  = 78;
  ram[4090]  = 79;
  ram[4091]  = 79;
  ram[4092]  = 78;
  ram[4093]  = 78;
  ram[4094]  = 77;
  ram[4095]  = 76;
end

always @(posedge clock) begin
  dout <= ram[address];
end

endmodule
