module rom_snaker (clock, address, q);
input clock;
output [7:0] q;
input [11:0] address;
reg [7:0] dout;
reg [7:0] ram [4095:0];
assign q = dout;

initial begin
  ram[0]  = 57;
  ram[1]  = 62;
  ram[2]  = 60;
  ram[3]  = 60;
  ram[4]  = 61;
  ram[5]  = 59;
  ram[6]  = 61;
  ram[7]  = 61;
  ram[8]  = 60;
  ram[9]  = 60;
  ram[10]  = 60;
  ram[11]  = 60;
  ram[12]  = 59;
  ram[13]  = 59;
  ram[14]  = 59;
  ram[15]  = 59;
  ram[16]  = 60;
  ram[17]  = 60;
  ram[18]  = 60;
  ram[19]  = 60;
  ram[20]  = 60;
  ram[21]  = 60;
  ram[22]  = 60;
  ram[23]  = 60;
  ram[24]  = 60;
  ram[25]  = 60;
  ram[26]  = 60;
  ram[27]  = 60;
  ram[28]  = 60;
  ram[29]  = 60;
  ram[30]  = 60;
  ram[31]  = 60;
  ram[32]  = 60;
  ram[33]  = 60;
  ram[34]  = 60;
  ram[35]  = 60;
  ram[36]  = 60;
  ram[37]  = 60;
  ram[38]  = 60;
  ram[39]  = 60;
  ram[40]  = 60;
  ram[41]  = 60;
  ram[42]  = 60;
  ram[43]  = 60;
  ram[44]  = 60;
  ram[45]  = 60;
  ram[46]  = 60;
  ram[47]  = 60;
  ram[48]  = 61;
  ram[49]  = 61;
  ram[50]  = 61;
  ram[51]  = 61;
  ram[52]  = 61;
  ram[53]  = 61;
  ram[54]  = 61;
  ram[55]  = 61;
  ram[56]  = 60;
  ram[57]  = 61;
  ram[58]  = 61;
  ram[59]  = 61;
  ram[60]  = 61;
  ram[61]  = 61;
  ram[62]  = 60;
  ram[63]  = 58;
  ram[64]  = 60;
  ram[65]  = 64;
  ram[66]  = 62;
  ram[67]  = 62;
  ram[68]  = 64;
  ram[69]  = 62;
  ram[70]  = 64;
  ram[71]  = 63;
  ram[72]  = 63;
  ram[73]  = 63;
  ram[74]  = 63;
  ram[75]  = 63;
  ram[76]  = 62;
  ram[77]  = 62;
  ram[78]  = 62;
  ram[79]  = 62;
  ram[80]  = 62;
  ram[81]  = 62;
  ram[82]  = 62;
  ram[83]  = 62;
  ram[84]  = 62;
  ram[85]  = 62;
  ram[86]  = 62;
  ram[87]  = 62;
  ram[88]  = 62;
  ram[89]  = 62;
  ram[90]  = 62;
  ram[91]  = 62;
  ram[92]  = 62;
  ram[93]  = 62;
  ram[94]  = 62;
  ram[95]  = 62;
  ram[96]  = 62;
  ram[97]  = 62;
  ram[98]  = 62;
  ram[99]  = 62;
  ram[100]  = 62;
  ram[101]  = 62;
  ram[102]  = 62;
  ram[103]  = 62;
  ram[104]  = 62;
  ram[105]  = 62;
  ram[106]  = 62;
  ram[107]  = 62;
  ram[108]  = 62;
  ram[109]  = 62;
  ram[110]  = 62;
  ram[111]  = 62;
  ram[112]  = 63;
  ram[113]  = 63;
  ram[114]  = 63;
  ram[115]  = 63;
  ram[116]  = 63;
  ram[117]  = 63;
  ram[118]  = 63;
  ram[119]  = 63;
  ram[120]  = 63;
  ram[121]  = 63;
  ram[122]  = 63;
  ram[123]  = 63;
  ram[124]  = 64;
  ram[125]  = 64;
  ram[126]  = 63;
  ram[127]  = 60;
  ram[128]  = 61;
  ram[129]  = 65;
  ram[130]  = 63;
  ram[131]  = 64;
  ram[132]  = 65;
  ram[133]  = 64;
  ram[134]  = 64;
  ram[135]  = 64;
  ram[136]  = 65;
  ram[137]  = 65;
  ram[138]  = 64;
  ram[139]  = 64;
  ram[140]  = 64;
  ram[141]  = 64;
  ram[142]  = 63;
  ram[143]  = 63;
  ram[144]  = 64;
  ram[145]  = 64;
  ram[146]  = 64;
  ram[147]  = 64;
  ram[148]  = 64;
  ram[149]  = 64;
  ram[150]  = 64;
  ram[151]  = 64;
  ram[152]  = 64;
  ram[153]  = 64;
  ram[154]  = 64;
  ram[155]  = 64;
  ram[156]  = 64;
  ram[157]  = 64;
  ram[158]  = 64;
  ram[159]  = 64;
  ram[160]  = 64;
  ram[161]  = 64;
  ram[162]  = 64;
  ram[163]  = 64;
  ram[164]  = 64;
  ram[165]  = 64;
  ram[166]  = 64;
  ram[167]  = 64;
  ram[168]  = 64;
  ram[169]  = 64;
  ram[170]  = 64;
  ram[171]  = 64;
  ram[172]  = 64;
  ram[173]  = 64;
  ram[174]  = 64;
  ram[175]  = 64;
  ram[176]  = 64;
  ram[177]  = 64;
  ram[178]  = 64;
  ram[179]  = 64;
  ram[180]  = 64;
  ram[181]  = 64;
  ram[182]  = 64;
  ram[183]  = 64;
  ram[184]  = 64;
  ram[185]  = 64;
  ram[186]  = 64;
  ram[187]  = 64;
  ram[188]  = 64;
  ram[189]  = 65;
  ram[190]  = 63;
  ram[191]  = 61;
  ram[192]  = 61;
  ram[193]  = 64;
  ram[194]  = 62;
  ram[195]  = 63;
  ram[196]  = 65;
  ram[197]  = 64;
  ram[198]  = 64;
  ram[199]  = 63;
  ram[200]  = 65;
  ram[201]  = 65;
  ram[202]  = 65;
  ram[203]  = 65;
  ram[204]  = 65;
  ram[205]  = 65;
  ram[206]  = 64;
  ram[207]  = 64;
  ram[208]  = 64;
  ram[209]  = 64;
  ram[210]  = 64;
  ram[211]  = 64;
  ram[212]  = 64;
  ram[213]  = 64;
  ram[214]  = 64;
  ram[215]  = 64;
  ram[216]  = 64;
  ram[217]  = 64;
  ram[218]  = 64;
  ram[219]  = 64;
  ram[220]  = 64;
  ram[221]  = 64;
  ram[222]  = 64;
  ram[223]  = 64;
  ram[224]  = 64;
  ram[225]  = 64;
  ram[226]  = 64;
  ram[227]  = 64;
  ram[228]  = 64;
  ram[229]  = 64;
  ram[230]  = 64;
  ram[231]  = 64;
  ram[232]  = 64;
  ram[233]  = 64;
  ram[234]  = 64;
  ram[235]  = 64;
  ram[236]  = 64;
  ram[237]  = 64;
  ram[238]  = 64;
  ram[239]  = 64;
  ram[240]  = 64;
  ram[241]  = 64;
  ram[242]  = 64;
  ram[243]  = 64;
  ram[244]  = 64;
  ram[245]  = 64;
  ram[246]  = 64;
  ram[247]  = 64;
  ram[248]  = 63;
  ram[249]  = 64;
  ram[250]  = 64;
  ram[251]  = 63;
  ram[252]  = 64;
  ram[253]  = 64;
  ram[254]  = 63;
  ram[255]  = 61;
  ram[256]  = 61;
  ram[257]  = 65;
  ram[258]  = 63;
  ram[259]  = 63;
  ram[260]  = 65;
  ram[261]  = 64;
  ram[262]  = 65;
  ram[263]  = 64;
  ram[264]  = 66;
  ram[265]  = 66;
  ram[266]  = 66;
  ram[267]  = 66;
  ram[268]  = 65;
  ram[269]  = 65;
  ram[270]  = 65;
  ram[271]  = 65;
  ram[272]  = 66;
  ram[273]  = 66;
  ram[274]  = 66;
  ram[275]  = 66;
  ram[276]  = 66;
  ram[277]  = 66;
  ram[278]  = 66;
  ram[279]  = 66;
  ram[280]  = 66;
  ram[281]  = 66;
  ram[282]  = 66;
  ram[283]  = 66;
  ram[284]  = 66;
  ram[285]  = 66;
  ram[286]  = 66;
  ram[287]  = 66;
  ram[288]  = 66;
  ram[289]  = 66;
  ram[290]  = 66;
  ram[291]  = 66;
  ram[292]  = 66;
  ram[293]  = 66;
  ram[294]  = 66;
  ram[295]  = 66;
  ram[296]  = 66;
  ram[297]  = 66;
  ram[298]  = 66;
  ram[299]  = 66;
  ram[300]  = 66;
  ram[301]  = 66;
  ram[302]  = 66;
  ram[303]  = 66;
  ram[304]  = 65;
  ram[305]  = 65;
  ram[306]  = 65;
  ram[307]  = 65;
  ram[308]  = 65;
  ram[309]  = 65;
  ram[310]  = 65;
  ram[311]  = 65;
  ram[312]  = 64;
  ram[313]  = 64;
  ram[314]  = 64;
  ram[315]  = 64;
  ram[316]  = 64;
  ram[317]  = 65;
  ram[318]  = 63;
  ram[319]  = 61;
  ram[320]  = 61;
  ram[321]  = 65;
  ram[322]  = 63;
  ram[323]  = 63;
  ram[324]  = 65;
  ram[325]  = 63;
  ram[326]  = 65;
  ram[327]  = 64;
  ram[328]  = 65;
  ram[329]  = 65;
  ram[330]  = 65;
  ram[331]  = 65;
  ram[332]  = 63;
  ram[333]  = 64;
  ram[334]  = 64;
  ram[335]  = 64;
  ram[336]  = 65;
  ram[337]  = 65;
  ram[338]  = 65;
  ram[339]  = 65;
  ram[340]  = 65;
  ram[341]  = 65;
  ram[342]  = 65;
  ram[343]  = 65;
  ram[344]  = 65;
  ram[345]  = 65;
  ram[346]  = 65;
  ram[347]  = 65;
  ram[348]  = 65;
  ram[349]  = 65;
  ram[350]  = 65;
  ram[351]  = 65;
  ram[352]  = 65;
  ram[353]  = 65;
  ram[354]  = 65;
  ram[355]  = 65;
  ram[356]  = 65;
  ram[357]  = 65;
  ram[358]  = 65;
  ram[359]  = 65;
  ram[360]  = 65;
  ram[361]  = 65;
  ram[362]  = 65;
  ram[363]  = 65;
  ram[364]  = 65;
  ram[365]  = 65;
  ram[366]  = 65;
  ram[367]  = 65;
  ram[368]  = 64;
  ram[369]  = 64;
  ram[370]  = 64;
  ram[371]  = 64;
  ram[372]  = 64;
  ram[373]  = 64;
  ram[374]  = 64;
  ram[375]  = 64;
  ram[376]  = 64;
  ram[377]  = 64;
  ram[378]  = 64;
  ram[379]  = 64;
  ram[380]  = 64;
  ram[381]  = 64;
  ram[382]  = 63;
  ram[383]  = 61;
  ram[384]  = 61;
  ram[385]  = 65;
  ram[386]  = 63;
  ram[387]  = 63;
  ram[388]  = 65;
  ram[389]  = 64;
  ram[390]  = 65;
  ram[391]  = 64;
  ram[392]  = 64;
  ram[393]  = 64;
  ram[394]  = 64;
  ram[395]  = 64;
  ram[396]  = 64;
  ram[397]  = 64;
  ram[398]  = 64;
  ram[399]  = 64;
  ram[400]  = 64;
  ram[401]  = 64;
  ram[402]  = 64;
  ram[403]  = 64;
  ram[404]  = 64;
  ram[405]  = 64;
  ram[406]  = 64;
  ram[407]  = 64;
  ram[408]  = 64;
  ram[409]  = 64;
  ram[410]  = 64;
  ram[411]  = 64;
  ram[412]  = 64;
  ram[413]  = 64;
  ram[414]  = 64;
  ram[415]  = 64;
  ram[416]  = 64;
  ram[417]  = 64;
  ram[418]  = 64;
  ram[419]  = 64;
  ram[420]  = 64;
  ram[421]  = 64;
  ram[422]  = 64;
  ram[423]  = 64;
  ram[424]  = 64;
  ram[425]  = 64;
  ram[426]  = 64;
  ram[427]  = 64;
  ram[428]  = 64;
  ram[429]  = 64;
  ram[430]  = 64;
  ram[431]  = 64;
  ram[432]  = 64;
  ram[433]  = 64;
  ram[434]  = 64;
  ram[435]  = 64;
  ram[436]  = 64;
  ram[437]  = 64;
  ram[438]  = 64;
  ram[439]  = 64;
  ram[440]  = 65;
  ram[441]  = 65;
  ram[442]  = 65;
  ram[443]  = 64;
  ram[444]  = 65;
  ram[445]  = 65;
  ram[446]  = 63;
  ram[447]  = 61;
  ram[448]  = 61;
  ram[449]  = 66;
  ram[450]  = 64;
  ram[451]  = 64;
  ram[452]  = 66;
  ram[453]  = 64;
  ram[454]  = 65;
  ram[455]  = 66;
  ram[456]  = 66;
  ram[457]  = 66;
  ram[458]  = 65;
  ram[459]  = 65;
  ram[460]  = 65;
  ram[461]  = 65;
  ram[462]  = 65;
  ram[463]  = 65;
  ram[464]  = 65;
  ram[465]  = 65;
  ram[466]  = 65;
  ram[467]  = 65;
  ram[468]  = 65;
  ram[469]  = 65;
  ram[470]  = 65;
  ram[471]  = 65;
  ram[472]  = 65;
  ram[473]  = 65;
  ram[474]  = 65;
  ram[475]  = 65;
  ram[476]  = 65;
  ram[477]  = 65;
  ram[478]  = 65;
  ram[479]  = 65;
  ram[480]  = 65;
  ram[481]  = 65;
  ram[482]  = 65;
  ram[483]  = 65;
  ram[484]  = 65;
  ram[485]  = 65;
  ram[486]  = 65;
  ram[487]  = 65;
  ram[488]  = 65;
  ram[489]  = 65;
  ram[490]  = 65;
  ram[491]  = 65;
  ram[492]  = 65;
  ram[493]  = 65;
  ram[494]  = 65;
  ram[495]  = 65;
  ram[496]  = 65;
  ram[497]  = 65;
  ram[498]  = 65;
  ram[499]  = 65;
  ram[500]  = 65;
  ram[501]  = 65;
  ram[502]  = 65;
  ram[503]  = 65;
  ram[504]  = 65;
  ram[505]  = 66;
  ram[506]  = 66;
  ram[507]  = 65;
  ram[508]  = 65;
  ram[509]  = 66;
  ram[510]  = 64;
  ram[511]  = 62;
  ram[512]  = 61;
  ram[513]  = 64;
  ram[514]  = 63;
  ram[515]  = 62;
  ram[516]  = 64;
  ram[517]  = 64;
  ram[518]  = 66;
  ram[519]  = 66;
  ram[520]  = 66;
  ram[521]  = 66;
  ram[522]  = 66;
  ram[523]  = 66;
  ram[524]  = 66;
  ram[525]  = 66;
  ram[526]  = 66;
  ram[527]  = 66;
  ram[528]  = 64;
  ram[529]  = 64;
  ram[530]  = 65;
  ram[531]  = 65;
  ram[532]  = 64;
  ram[533]  = 64;
  ram[534]  = 64;
  ram[535]  = 65;
  ram[536]  = 64;
  ram[537]  = 64;
  ram[538]  = 64;
  ram[539]  = 64;
  ram[540]  = 64;
  ram[541]  = 64;
  ram[542]  = 64;
  ram[543]  = 64;
  ram[544]  = 64;
  ram[545]  = 64;
  ram[546]  = 64;
  ram[547]  = 64;
  ram[548]  = 64;
  ram[549]  = 64;
  ram[550]  = 64;
  ram[551]  = 64;
  ram[552]  = 63;
  ram[553]  = 64;
  ram[554]  = 64;
  ram[555]  = 64;
  ram[556]  = 64;
  ram[557]  = 64;
  ram[558]  = 64;
  ram[559]  = 64;
  ram[560]  = 64;
  ram[561]  = 64;
  ram[562]  = 64;
  ram[563]  = 64;
  ram[564]  = 64;
  ram[565]  = 64;
  ram[566]  = 64;
  ram[567]  = 63;
  ram[568]  = 63;
  ram[569]  = 64;
  ram[570]  = 64;
  ram[571]  = 64;
  ram[572]  = 64;
  ram[573]  = 65;
  ram[574]  = 63;
  ram[575]  = 62;
  ram[576]  = 62;
  ram[577]  = 65;
  ram[578]  = 65;
  ram[579]  = 64;
  ram[580]  = 66;
  ram[581]  = 66;
  ram[582]  = 67;
  ram[583]  = 67;
  ram[584]  = 67;
  ram[585]  = 67;
  ram[586]  = 67;
  ram[587]  = 67;
  ram[588]  = 67;
  ram[589]  = 67;
  ram[590]  = 67;
  ram[591]  = 67;
  ram[592]  = 65;
  ram[593]  = 66;
  ram[594]  = 66;
  ram[595]  = 66;
  ram[596]  = 65;
  ram[597]  = 65;
  ram[598]  = 65;
  ram[599]  = 65;
  ram[600]  = 66;
  ram[601]  = 66;
  ram[602]  = 66;
  ram[603]  = 66;
  ram[604]  = 66;
  ram[605]  = 66;
  ram[606]  = 66;
  ram[607]  = 65;
  ram[608]  = 66;
  ram[609]  = 66;
  ram[610]  = 66;
  ram[611]  = 66;
  ram[612]  = 66;
  ram[613]  = 67;
  ram[614]  = 67;
  ram[615]  = 67;
  ram[616]  = 67;
  ram[617]  = 67;
  ram[618]  = 67;
  ram[619]  = 67;
  ram[620]  = 67;
  ram[621]  = 67;
  ram[622]  = 67;
  ram[623]  = 67;
  ram[624]  = 66;
  ram[625]  = 66;
  ram[626]  = 66;
  ram[627]  = 66;
  ram[628]  = 66;
  ram[629]  = 66;
  ram[630]  = 66;
  ram[631]  = 65;
  ram[632]  = 65;
  ram[633]  = 66;
  ram[634]  = 66;
  ram[635]  = 65;
  ram[636]  = 65;
  ram[637]  = 65;
  ram[638]  = 64;
  ram[639]  = 62;
  ram[640]  = 63;
  ram[641]  = 66;
  ram[642]  = 66;
  ram[643]  = 65;
  ram[644]  = 66;
  ram[645]  = 66;
  ram[646]  = 67;
  ram[647]  = 67;
  ram[648]  = 67;
  ram[649]  = 67;
  ram[650]  = 68;
  ram[651]  = 68;
  ram[652]  = 67;
  ram[653]  = 67;
  ram[654]  = 67;
  ram[655]  = 67;
  ram[656]  = 66;
  ram[657]  = 66;
  ram[658]  = 65;
  ram[659]  = 65;
  ram[660]  = 65;
  ram[661]  = 65;
  ram[662]  = 65;
  ram[663]  = 65;
  ram[664]  = 65;
  ram[665]  = 65;
  ram[666]  = 65;
  ram[667]  = 65;
  ram[668]  = 65;
  ram[669]  = 65;
  ram[670]  = 65;
  ram[671]  = 65;
  ram[672]  = 65;
  ram[673]  = 65;
  ram[674]  = 65;
  ram[675]  = 64;
  ram[676]  = 64;
  ram[677]  = 64;
  ram[678]  = 64;
  ram[679]  = 64;
  ram[680]  = 64;
  ram[681]  = 64;
  ram[682]  = 64;
  ram[683]  = 64;
  ram[684]  = 64;
  ram[685]  = 64;
  ram[686]  = 64;
  ram[687]  = 64;
  ram[688]  = 67;
  ram[689]  = 67;
  ram[690]  = 67;
  ram[691]  = 68;
  ram[692]  = 67;
  ram[693]  = 67;
  ram[694]  = 67;
  ram[695]  = 67;
  ram[696]  = 67;
  ram[697]  = 68;
  ram[698]  = 68;
  ram[699]  = 67;
  ram[700]  = 67;
  ram[701]  = 67;
  ram[702]  = 66;
  ram[703]  = 64;
  ram[704]  = 62;
  ram[705]  = 65;
  ram[706]  = 65;
  ram[707]  = 64;
  ram[708]  = 65;
  ram[709]  = 65;
  ram[710]  = 65;
  ram[711]  = 66;
  ram[712]  = 66;
  ram[713]  = 66;
  ram[714]  = 67;
  ram[715]  = 67;
  ram[716]  = 66;
  ram[717]  = 66;
  ram[718]  = 66;
  ram[719]  = 66;
  ram[720]  = 67;
  ram[721]  = 65;
  ram[722]  = 66;
  ram[723]  = 64;
  ram[724]  = 66;
  ram[725]  = 64;
  ram[726]  = 66;
  ram[727]  = 63;
  ram[728]  = 64;
  ram[729]  = 63;
  ram[730]  = 65;
  ram[731]  = 63;
  ram[732]  = 65;
  ram[733]  = 64;
  ram[734]  = 66;
  ram[735]  = 64;
  ram[736]  = 69;
  ram[737]  = 67;
  ram[738]  = 69;
  ram[739]  = 66;
  ram[740]  = 68;
  ram[741]  = 66;
  ram[742]  = 68;
  ram[743]  = 66;
  ram[744]  = 67;
  ram[745]  = 65;
  ram[746]  = 67;
  ram[747]  = 65;
  ram[748]  = 68;
  ram[749]  = 66;
  ram[750]  = 68;
  ram[751]  = 68;
  ram[752]  = 66;
  ram[753]  = 66;
  ram[754]  = 66;
  ram[755]  = 66;
  ram[756]  = 66;
  ram[757]  = 66;
  ram[758]  = 66;
  ram[759]  = 66;
  ram[760]  = 65;
  ram[761]  = 66;
  ram[762]  = 66;
  ram[763]  = 66;
  ram[764]  = 66;
  ram[765]  = 66;
  ram[766]  = 65;
  ram[767]  = 64;
  ram[768]  = 62;
  ram[769]  = 64;
  ram[770]  = 65;
  ram[771]  = 63;
  ram[772]  = 66;
  ram[773]  = 66;
  ram[774]  = 65;
  ram[775]  = 66;
  ram[776]  = 67;
  ram[777]  = 67;
  ram[778]  = 67;
  ram[779]  = 67;
  ram[780]  = 67;
  ram[781]  = 67;
  ram[782]  = 67;
  ram[783]  = 67;
  ram[784]  = 68;
  ram[785]  = 66;
  ram[786]  = 66;
  ram[787]  = 65;
  ram[788]  = 67;
  ram[789]  = 66;
  ram[790]  = 66;
  ram[791]  = 64;
  ram[792]  = 66;
  ram[793]  = 65;
  ram[794]  = 66;
  ram[795]  = 66;
  ram[796]  = 67;
  ram[797]  = 66;
  ram[798]  = 67;
  ram[799]  = 66;
  ram[800]  = 65;
  ram[801]  = 65;
  ram[802]  = 66;
  ram[803]  = 65;
  ram[804]  = 66;
  ram[805]  = 65;
  ram[806]  = 66;
  ram[807]  = 65;
  ram[808]  = 66;
  ram[809]  = 65;
  ram[810]  = 66;
  ram[811]  = 65;
  ram[812]  = 66;
  ram[813]  = 65;
  ram[814]  = 66;
  ram[815]  = 65;
  ram[816]  = 66;
  ram[817]  = 67;
  ram[818]  = 67;
  ram[819]  = 67;
  ram[820]  = 67;
  ram[821]  = 67;
  ram[822]  = 67;
  ram[823]  = 67;
  ram[824]  = 65;
  ram[825]  = 66;
  ram[826]  = 66;
  ram[827]  = 65;
  ram[828]  = 65;
  ram[829]  = 66;
  ram[830]  = 65;
  ram[831]  = 64;
  ram[832]  = 62;
  ram[833]  = 64;
  ram[834]  = 65;
  ram[835]  = 64;
  ram[836]  = 67;
  ram[837]  = 67;
  ram[838]  = 66;
  ram[839]  = 66;
  ram[840]  = 67;
  ram[841]  = 67;
  ram[842]  = 67;
  ram[843]  = 67;
  ram[844]  = 67;
  ram[845]  = 67;
  ram[846]  = 67;
  ram[847]  = 67;
  ram[848]  = 67;
  ram[849]  = 67;
  ram[850]  = 69;
  ram[851]  = 67;
  ram[852]  = 69;
  ram[853]  = 67;
  ram[854]  = 69;
  ram[855]  = 67;
  ram[856]  = 70;
  ram[857]  = 68;
  ram[858]  = 69;
  ram[859]  = 67;
  ram[860]  = 69;
  ram[861]  = 67;
  ram[862]  = 68;
  ram[863]  = 66;
  ram[864]  = 70;
  ram[865]  = 68;
  ram[866]  = 70;
  ram[867]  = 69;
  ram[868]  = 71;
  ram[869]  = 70;
  ram[870]  = 72;
  ram[871]  = 71;
  ram[872]  = 72;
  ram[873]  = 70;
  ram[874]  = 72;
  ram[875]  = 70;
  ram[876]  = 72;
  ram[877]  = 70;
  ram[878]  = 72;
  ram[879]  = 70;
  ram[880]  = 67;
  ram[881]  = 67;
  ram[882]  = 67;
  ram[883]  = 67;
  ram[884]  = 67;
  ram[885]  = 67;
  ram[886]  = 67;
  ram[887]  = 67;
  ram[888]  = 67;
  ram[889]  = 67;
  ram[890]  = 67;
  ram[891]  = 66;
  ram[892]  = 65;
  ram[893]  = 65;
  ram[894]  = 65;
  ram[895]  = 63;
  ram[896]  = 60;
  ram[897]  = 63;
  ram[898]  = 64;
  ram[899]  = 63;
  ram[900]  = 66;
  ram[901]  = 66;
  ram[902]  = 66;
  ram[903]  = 67;
  ram[904]  = 67;
  ram[905]  = 67;
  ram[906]  = 67;
  ram[907]  = 67;
  ram[908]  = 66;
  ram[909]  = 66;
  ram[910]  = 66;
  ram[911]  = 66;
  ram[912]  = 68;
  ram[913]  = 68;
  ram[914]  = 69;
  ram[915]  = 68;
  ram[916]  = 69;
  ram[917]  = 68;
  ram[918]  = 69;
  ram[919]  = 69;
  ram[920]  = 69;
  ram[921]  = 68;
  ram[922]  = 69;
  ram[923]  = 68;
  ram[924]  = 69;
  ram[925]  = 68;
  ram[926]  = 69;
  ram[927]  = 68;
  ram[928]  = 69;
  ram[929]  = 68;
  ram[930]  = 69;
  ram[931]  = 68;
  ram[932]  = 69;
  ram[933]  = 68;
  ram[934]  = 69;
  ram[935]  = 68;
  ram[936]  = 69;
  ram[937]  = 68;
  ram[938]  = 69;
  ram[939]  = 68;
  ram[940]  = 69;
  ram[941]  = 68;
  ram[942]  = 69;
  ram[943]  = 68;
  ram[944]  = 67;
  ram[945]  = 66;
  ram[946]  = 66;
  ram[947]  = 66;
  ram[948]  = 66;
  ram[949]  = 66;
  ram[950]  = 66;
  ram[951]  = 66;
  ram[952]  = 66;
  ram[953]  = 67;
  ram[954]  = 66;
  ram[955]  = 65;
  ram[956]  = 65;
  ram[957]  = 65;
  ram[958]  = 64;
  ram[959]  = 63;
  ram[960]  = 58;
  ram[961]  = 61;
  ram[962]  = 62;
  ram[963]  = 61;
  ram[964]  = 64;
  ram[965]  = 66;
  ram[966]  = 65;
  ram[967]  = 68;
  ram[968]  = 67;
  ram[969]  = 67;
  ram[970]  = 67;
  ram[971]  = 67;
  ram[972]  = 67;
  ram[973]  = 67;
  ram[974]  = 67;
  ram[975]  = 67;
  ram[976]  = 67;
  ram[977]  = 68;
  ram[978]  = 67;
  ram[979]  = 67;
  ram[980]  = 67;
  ram[981]  = 67;
  ram[982]  = 68;
  ram[983]  = 69;
  ram[984]  = 67;
  ram[985]  = 68;
  ram[986]  = 68;
  ram[987]  = 68;
  ram[988]  = 69;
  ram[989]  = 70;
  ram[990]  = 71;
  ram[991]  = 70;
  ram[992]  = 71;
  ram[993]  = 71;
  ram[994]  = 70;
  ram[995]  = 69;
  ram[996]  = 68;
  ram[997]  = 68;
  ram[998]  = 68;
  ram[999]  = 68;
  ram[1000]  = 68;
  ram[1001]  = 68;
  ram[1002]  = 67;
  ram[1003]  = 67;
  ram[1004]  = 69;
  ram[1005]  = 69;
  ram[1006]  = 70;
  ram[1007]  = 69;
  ram[1008]  = 68;
  ram[1009]  = 66;
  ram[1010]  = 68;
  ram[1011]  = 69;
  ram[1012]  = 67;
  ram[1013]  = 67;
  ram[1014]  = 67;
  ram[1015]  = 67;
  ram[1016]  = 67;
  ram[1017]  = 67;
  ram[1018]  = 65;
  ram[1019]  = 64;
  ram[1020]  = 63;
  ram[1021]  = 64;
  ram[1022]  = 64;
  ram[1023]  = 62;
  ram[1024]  = 57;
  ram[1025]  = 62;
  ram[1026]  = 63;
  ram[1027]  = 59;
  ram[1028]  = 64;
  ram[1029]  = 62;
  ram[1030]  = 65;
  ram[1031]  = 46;
  ram[1032]  = 50;
  ram[1033]  = 55;
  ram[1034]  = 53;
  ram[1035]  = 50;
  ram[1036]  = 54;
  ram[1037]  = 47;
  ram[1038]  = 63;
  ram[1039]  = 65;
  ram[1040]  = 57;
  ram[1041]  = 50;
  ram[1042]  = 63;
  ram[1043]  = 62;
  ram[1044]  = 65;
  ram[1045]  = 62;
  ram[1046]  = 64;
  ram[1047]  = 61;
  ram[1048]  = 51;
  ram[1049]  = 59;
  ram[1050]  = 63;
  ram[1051]  = 67;
  ram[1052]  = 65;
  ram[1053]  = 59;
  ram[1054]  = 48;
  ram[1055]  = 53;
  ram[1056]  = 53;
  ram[1057]  = 50;
  ram[1058]  = 50;
  ram[1059]  = 65;
  ram[1060]  = 67;
  ram[1061]  = 66;
  ram[1062]  = 61;
  ram[1063]  = 52;
  ram[1064]  = 58;
  ram[1065]  = 64;
  ram[1066]  = 62;
  ram[1067]  = 62;
  ram[1068]  = 61;
  ram[1069]  = 67;
  ram[1070]  = 54;
  ram[1071]  = 53;
  ram[1072]  = 66;
  ram[1073]  = 64;
  ram[1074]  = 49;
  ram[1075]  = 60;
  ram[1076]  = 48;
  ram[1077]  = 54;
  ram[1078]  = 50;
  ram[1079]  = 52;
  ram[1080]  = 54;
  ram[1081]  = 58;
  ram[1082]  = 49;
  ram[1083]  = 58;
  ram[1084]  = 66;
  ram[1085]  = 62;
  ram[1086]  = 61;
  ram[1087]  = 61;
  ram[1088]  = 58;
  ram[1089]  = 65;
  ram[1090]  = 59;
  ram[1091]  = 62;
  ram[1092]  = 71;
  ram[1093]  = 57;
  ram[1094]  = 69;
  ram[1095]  = 135;
  ram[1096]  = 118;
  ram[1097]  = 118;
  ram[1098]  = 115;
  ram[1099]  = 129;
  ram[1100]  = 111;
  ram[1101]  = 142;
  ram[1102]  = 68;
  ram[1103]  = 45;
  ram[1104]  = 123;
  ram[1105]  = 129;
  ram[1106]  = 51;
  ram[1107]  = 66;
  ram[1108]  = 59;
  ram[1109]  = 64;
  ram[1110]  = 65;
  ram[1111]  = 80;
  ram[1112]  = 136;
  ram[1113]  = 96;
  ram[1114]  = 59;
  ram[1115]  = 67;
  ram[1116]  = 52;
  ram[1117]  = 107;
  ram[1118]  = 130;
  ram[1119]  = 120;
  ram[1120]  = 121;
  ram[1121]  = 121;
  ram[1122]  = 111;
  ram[1123]  = 59;
  ram[1124]  = 63;
  ram[1125]  = 57;
  ram[1126]  = 82;
  ram[1127]  = 137;
  ram[1128]  = 90;
  ram[1129]  = 57;
  ram[1130]  = 65;
  ram[1131]  = 57;
  ram[1132]  = 68;
  ram[1133]  = 56;
  ram[1134]  = 130;
  ram[1135]  = 144;
  ram[1136]  = 50;
  ram[1137]  = 56;
  ram[1138]  = 137;
  ram[1139]  = 117;
  ram[1140]  = 125;
  ram[1141]  = 112;
  ram[1142]  = 125;
  ram[1143]  = 117;
  ram[1144]  = 125;
  ram[1145]  = 117;
  ram[1146]  = 131;
  ram[1147]  = 79;
  ram[1148]  = 57;
  ram[1149]  = 61;
  ram[1150]  = 68;
  ram[1151]  = 65;
  ram[1152]  = 72;
  ram[1153]  = 61;
  ram[1154]  = 76;
  ram[1155]  = 66;
  ram[1156]  = 61;
  ram[1157]  = 46;
  ram[1158]  = 82;
  ram[1159]  = 204;
  ram[1160]  = 196;
  ram[1161]  = 203;
  ram[1162]  = 201;
  ram[1163]  = 201;
  ram[1164]  = 201;
  ram[1165]  = 203;
  ram[1166]  = 76;
  ram[1167]  = 28;
  ram[1168]  = 196;
  ram[1169]  = 194;
  ram[1170]  = 44;
  ram[1171]  = 61;
  ram[1172]  = 66;
  ram[1173]  = 61;
  ram[1174]  = 61;
  ram[1175]  = 103;
  ram[1176]  = 198;
  ram[1177]  = 132;
  ram[1178]  = 46;
  ram[1179]  = 48;
  ram[1180]  = 38;
  ram[1181]  = 165;
  ram[1182]  = 201;
  ram[1183]  = 199;
  ram[1184]  = 200;
  ram[1185]  = 195;
  ram[1186]  = 177;
  ram[1187]  = 29;
  ram[1188]  = 41;
  ram[1189]  = 53;
  ram[1190]  = 105;
  ram[1191]  = 200;
  ram[1192]  = 111;
  ram[1193]  = 52;
  ram[1194]  = 54;
  ram[1195]  = 67;
  ram[1196]  = 40;
  ram[1197]  = 15;
  ram[1198]  = 211;
  ram[1199]  = 215;
  ram[1200]  = 22;
  ram[1201]  = 47;
  ram[1202]  = 196;
  ram[1203]  = 185;
  ram[1204]  = 198;
  ram[1205]  = 193;
  ram[1206]  = 197;
  ram[1207]  = 192;
  ram[1208]  = 196;
  ram[1209]  = 195;
  ram[1210]  = 201;
  ram[1211]  = 93;
  ram[1212]  = 54;
  ram[1213]  = 64;
  ram[1214]  = 66;
  ram[1215]  = 62;
  ram[1216]  = 64;
  ram[1217]  = 69;
  ram[1218]  = 75;
  ram[1219]  = 67;
  ram[1220]  = 73;
  ram[1221]  = 158;
  ram[1222]  = 125;
  ram[1223]  = 84;
  ram[1224]  = 86;
  ram[1225]  = 87;
  ram[1226]  = 82;
  ram[1227]  = 89;
  ram[1228]  = 87;
  ram[1229]  = 99;
  ram[1230]  = 60;
  ram[1231]  = 31;
  ram[1232]  = 183;
  ram[1233]  = 187;
  ram[1234]  = 38;
  ram[1235]  = 60;
  ram[1236]  = 67;
  ram[1237]  = 69;
  ram[1238]  = 57;
  ram[1239]  = 94;
  ram[1240]  = 198;
  ram[1241]  = 107;
  ram[1242]  = 33;
  ram[1243]  = 113;
  ram[1244]  = 154;
  ram[1245]  = 86;
  ram[1246]  = 86;
  ram[1247]  = 87;
  ram[1248]  = 87;
  ram[1249]  = 80;
  ram[1250]  = 81;
  ram[1251]  = 157;
  ram[1252]  = 125;
  ram[1253]  = 38;
  ram[1254]  = 88;
  ram[1255]  = 189;
  ram[1256]  = 102;
  ram[1257]  = 52;
  ram[1258]  = 59;
  ram[1259]  = 47;
  ram[1260]  = 135;
  ram[1261]  = 162;
  ram[1262]  = 84;
  ram[1263]  = 94;
  ram[1264]  = 46;
  ram[1265]  = 49;
  ram[1266]  = 196;
  ram[1267]  = 148;
  ram[1268]  = 67;
  ram[1269]  = 78;
  ram[1270]  = 90;
  ram[1271]  = 80;
  ram[1272]  = 89;
  ram[1273]  = 88;
  ram[1274]  = 94;
  ram[1275]  = 62;
  ram[1276]  = 61;
  ram[1277]  = 62;
  ram[1278]  = 59;
  ram[1279]  = 64;
  ram[1280]  = 63;
  ram[1281]  = 68;
  ram[1282]  = 63;
  ram[1283]  = 60;
  ram[1284]  = 69;
  ram[1285]  = 192;
  ram[1286]  = 168;
  ram[1287]  = 24;
  ram[1288]  = 51;
  ram[1289]  = 52;
  ram[1290]  = 54;
  ram[1291]  = 45;
  ram[1292]  = 55;
  ram[1293]  = 52;
  ram[1294]  = 57;
  ram[1295]  = 28;
  ram[1296]  = 189;
  ram[1297]  = 191;
  ram[1298]  = 11;
  ram[1299]  = 37;
  ram[1300]  = 68;
  ram[1301]  = 66;
  ram[1302]  = 65;
  ram[1303]  = 91;
  ram[1304]  = 192;
  ram[1305]  = 124;
  ram[1306]  = 26;
  ram[1307]  = 134;
  ram[1308]  = 196;
  ram[1309]  = 76;
  ram[1310]  = 41;
  ram[1311]  = 51;
  ram[1312]  = 57;
  ram[1313]  = 47;
  ram[1314]  = 66;
  ram[1315]  = 191;
  ram[1316]  = 158;
  ram[1317]  = 34;
  ram[1318]  = 98;
  ram[1319]  = 196;
  ram[1320]  = 101;
  ram[1321]  = 51;
  ram[1322]  = 46;
  ram[1323]  = 16;
  ram[1324]  = 203;
  ram[1325]  = 212;
  ram[1326]  = 44;
  ram[1327]  = 55;
  ram[1328]  = 58;
  ram[1329]  = 51;
  ram[1330]  = 201;
  ram[1331]  = 161;
  ram[1332]  = 23;
  ram[1333]  = 48;
  ram[1334]  = 49;
  ram[1335]  = 52;
  ram[1336]  = 57;
  ram[1337]  = 59;
  ram[1338]  = 59;
  ram[1339]  = 60;
  ram[1340]  = 62;
  ram[1341]  = 59;
  ram[1342]  = 66;
  ram[1343]  = 63;
  ram[1344]  = 62;
  ram[1345]  = 68;
  ram[1346]  = 63;
  ram[1347]  = 62;
  ram[1348]  = 57;
  ram[1349]  = 189;
  ram[1350]  = 137;
  ram[1351]  = 47;
  ram[1352]  = 61;
  ram[1353]  = 61;
  ram[1354]  = 65;
  ram[1355]  = 59;
  ram[1356]  = 54;
  ram[1357]  = 67;
  ram[1358]  = 62;
  ram[1359]  = 27;
  ram[1360]  = 177;
  ram[1361]  = 167;
  ram[1362]  = 154;
  ram[1363]  = 166;
  ram[1364]  = 39;
  ram[1365]  = 59;
  ram[1366]  = 55;
  ram[1367]  = 94;
  ram[1368]  = 194;
  ram[1369]  = 103;
  ram[1370]  = 26;
  ram[1371]  = 122;
  ram[1372]  = 179;
  ram[1373]  = 76;
  ram[1374]  = 54;
  ram[1375]  = 65;
  ram[1376]  = 63;
  ram[1377]  = 65;
  ram[1378]  = 72;
  ram[1379]  = 183;
  ram[1380]  = 144;
  ram[1381]  = 30;
  ram[1382]  = 90;
  ram[1383]  = 190;
  ram[1384]  = 94;
  ram[1385]  = 36;
  ram[1386]  = 142;
  ram[1387]  = 196;
  ram[1388]  = 73;
  ram[1389]  = 72;
  ram[1390]  = 59;
  ram[1391]  = 59;
  ram[1392]  = 64;
  ram[1393]  = 37;
  ram[1394]  = 197;
  ram[1395]  = 158;
  ram[1396]  = 32;
  ram[1397]  = 67;
  ram[1398]  = 65;
  ram[1399]  = 62;
  ram[1400]  = 63;
  ram[1401]  = 67;
  ram[1402]  = 67;
  ram[1403]  = 64;
  ram[1404]  = 66;
  ram[1405]  = 57;
  ram[1406]  = 61;
  ram[1407]  = 58;
  ram[1408]  = 63;
  ram[1409]  = 67;
  ram[1410]  = 63;
  ram[1411]  = 62;
  ram[1412]  = 66;
  ram[1413]  = 191;
  ram[1414]  = 139;
  ram[1415]  = 0;
  ram[1416]  = 35;
  ram[1417]  = 35;
  ram[1418]  = 31;
  ram[1419]  = 37;
  ram[1420]  = 52;
  ram[1421]  = 62;
  ram[1422]  = 64;
  ram[1423]  = 31;
  ram[1424]  = 184;
  ram[1425]  = 177;
  ram[1426]  = 197;
  ram[1427]  = 194;
  ram[1428]  = 4;
  ram[1429]  = 41;
  ram[1430]  = 45;
  ram[1431]  = 95;
  ram[1432]  = 198;
  ram[1433]  = 115;
  ram[1434]  = 23;
  ram[1435]  = 130;
  ram[1436]  = 185;
  ram[1437]  = 51;
  ram[1438]  = 15;
  ram[1439]  = 29;
  ram[1440]  = 32;
  ram[1441]  = 17;
  ram[1442]  = 50;
  ram[1443]  = 186;
  ram[1444]  = 150;
  ram[1445]  = 29;
  ram[1446]  = 96;
  ram[1447]  = 203;
  ram[1448]  = 89;
  ram[1449]  = 0;
  ram[1450]  = 171;
  ram[1451]  = 225;
  ram[1452]  = 66;
  ram[1453]  = 53;
  ram[1454]  = 60;
  ram[1455]  = 68;
  ram[1456]  = 59;
  ram[1457]  = 56;
  ram[1458]  = 200;
  ram[1459]  = 151;
  ram[1460]  = 0;
  ram[1461]  = 34;
  ram[1462]  = 33;
  ram[1463]  = 32;
  ram[1464]  = 38;
  ram[1465]  = 52;
  ram[1466]  = 64;
  ram[1467]  = 64;
  ram[1468]  = 64;
  ram[1469]  = 61;
  ram[1470]  = 66;
  ram[1471]  = 65;
  ram[1472]  = 64;
  ram[1473]  = 63;
  ram[1474]  = 71;
  ram[1475]  = 60;
  ram[1476]  = 67;
  ram[1477]  = 181;
  ram[1478]  = 164;
  ram[1479]  = 188;
  ram[1480]  = 177;
  ram[1481]  = 194;
  ram[1482]  = 186;
  ram[1483]  = 202;
  ram[1484]  = 96;
  ram[1485]  = 57;
  ram[1486]  = 63;
  ram[1487]  = 29;
  ram[1488]  = 186;
  ram[1489]  = 189;
  ram[1490]  = 1;
  ram[1491]  = 22;
  ram[1492]  = 202;
  ram[1493]  = 170;
  ram[1494]  = 33;
  ram[1495]  = 85;
  ram[1496]  = 199;
  ram[1497]  = 110;
  ram[1498]  = 14;
  ram[1499]  = 124;
  ram[1500]  = 173;
  ram[1501]  = 169;
  ram[1502]  = 193;
  ram[1503]  = 187;
  ram[1504]  = 184;
  ram[1505]  = 189;
  ram[1506]  = 168;
  ram[1507]  = 174;
  ram[1508]  = 140;
  ram[1509]  = 23;
  ram[1510]  = 98;
  ram[1511]  = 184;
  ram[1512]  = 165;
  ram[1513]  = 215;
  ram[1514]  = 72;
  ram[1515]  = 43;
  ram[1516]  = 54;
  ram[1517]  = 63;
  ram[1518]  = 62;
  ram[1519]  = 53;
  ram[1520]  = 60;
  ram[1521]  = 49;
  ram[1522]  = 195;
  ram[1523]  = 163;
  ram[1524]  = 189;
  ram[1525]  = 179;
  ram[1526]  = 188;
  ram[1527]  = 186;
  ram[1528]  = 199;
  ram[1529]  = 112;
  ram[1530]  = 57;
  ram[1531]  = 66;
  ram[1532]  = 63;
  ram[1533]  = 59;
  ram[1534]  = 63;
  ram[1535]  = 57;
  ram[1536]  = 64;
  ram[1537]  = 68;
  ram[1538]  = 69;
  ram[1539]  = 65;
  ram[1540]  = 75;
  ram[1541]  = 199;
  ram[1542]  = 197;
  ram[1543]  = 201;
  ram[1544]  = 200;
  ram[1545]  = 203;
  ram[1546]  = 201;
  ram[1547]  = 212;
  ram[1548]  = 79;
  ram[1549]  = 28;
  ram[1550]  = 63;
  ram[1551]  = 31;
  ram[1552]  = 196;
  ram[1553]  = 200;
  ram[1554]  = 20;
  ram[1555]  = 54;
  ram[1556]  = 216;
  ram[1557]  = 172;
  ram[1558]  = 2;
  ram[1559]  = 73;
  ram[1560]  = 197;
  ram[1561]  = 125;
  ram[1562]  = 28;
  ram[1563]  = 131;
  ram[1564]  = 177;
  ram[1565]  = 189;
  ram[1566]  = 196;
  ram[1567]  = 204;
  ram[1568]  = 198;
  ram[1569]  = 196;
  ram[1570]  = 186;
  ram[1571]  = 178;
  ram[1572]  = 144;
  ram[1573]  = 30;
  ram[1574]  = 93;
  ram[1575]  = 185;
  ram[1576]  = 186;
  ram[1577]  = 219;
  ram[1578]  = 69;
  ram[1579]  = 25;
  ram[1580]  = 58;
  ram[1581]  = 63;
  ram[1582]  = 55;
  ram[1583]  = 60;
  ram[1584]  = 58;
  ram[1585]  = 51;
  ram[1586]  = 198;
  ram[1587]  = 175;
  ram[1588]  = 202;
  ram[1589]  = 196;
  ram[1590]  = 203;
  ram[1591]  = 197;
  ram[1592]  = 204;
  ram[1593]  = 105;
  ram[1594]  = 59;
  ram[1595]  = 64;
  ram[1596]  = 67;
  ram[1597]  = 65;
  ram[1598]  = 61;
  ram[1599]  = 62;
  ram[1600]  = 66;
  ram[1601]  = 61;
  ram[1602]  = 66;
  ram[1603]  = 64;
  ram[1604]  = 67;
  ram[1605]  = 37;
  ram[1606]  = 29;
  ram[1607]  = 35;
  ram[1608]  = 25;
  ram[1609]  = 34;
  ram[1610]  = 26;
  ram[1611]  = 7;
  ram[1612]  = 147;
  ram[1613]  = 223;
  ram[1614]  = 81;
  ram[1615]  = 22;
  ram[1616]  = 195;
  ram[1617]  = 206;
  ram[1618]  = 38;
  ram[1619]  = 57;
  ram[1620]  = 24;
  ram[1621]  = 56;
  ram[1622]  = 215;
  ram[1623]  = 191;
  ram[1624]  = 185;
  ram[1625]  = 119;
  ram[1626]  = 19;
  ram[1627]  = 130;
  ram[1628]  = 186;
  ram[1629]  = 54;
  ram[1630]  = 24;
  ram[1631]  = 27;
  ram[1632]  = 24;
  ram[1633]  = 22;
  ram[1634]  = 39;
  ram[1635]  = 181;
  ram[1636]  = 146;
  ram[1637]  = 28;
  ram[1638]  = 91;
  ram[1639]  = 201;
  ram[1640]  = 82;
  ram[1641]  = 0;
  ram[1642]  = 158;
  ram[1643]  = 226;
  ram[1644]  = 81;
  ram[1645]  = 48;
  ram[1646]  = 60;
  ram[1647]  = 57;
  ram[1648]  = 60;
  ram[1649]  = 47;
  ram[1650]  = 206;
  ram[1651]  = 148;
  ram[1652]  = 0;
  ram[1653]  = 26;
  ram[1654]  = 28;
  ram[1655]  = 28;
  ram[1656]  = 39;
  ram[1657]  = 58;
  ram[1658]  = 64;
  ram[1659]  = 66;
  ram[1660]  = 63;
  ram[1661]  = 58;
  ram[1662]  = 65;
  ram[1663]  = 60;
  ram[1664]  = 60;
  ram[1665]  = 62;
  ram[1666]  = 68;
  ram[1667]  = 65;
  ram[1668]  = 55;
  ram[1669]  = 61;
  ram[1670]  = 59;
  ram[1671]  = 60;
  ram[1672]  = 66;
  ram[1673]  = 64;
  ram[1674]  = 62;
  ram[1675]  = 42;
  ram[1676]  = 143;
  ram[1677]  = 209;
  ram[1678]  = 63;
  ram[1679]  = 20;
  ram[1680]  = 195;
  ram[1681]  = 196;
  ram[1682]  = 39;
  ram[1683]  = 57;
  ram[1684]  = 51;
  ram[1685]  = 84;
  ram[1686]  = 204;
  ram[1687]  = 182;
  ram[1688]  = 188;
  ram[1689]  = 114;
  ram[1690]  = 24;
  ram[1691]  = 135;
  ram[1692]  = 192;
  ram[1693]  = 74;
  ram[1694]  = 56;
  ram[1695]  = 60;
  ram[1696]  = 61;
  ram[1697]  = 53;
  ram[1698]  = 58;
  ram[1699]  = 198;
  ram[1700]  = 147;
  ram[1701]  = 21;
  ram[1702]  = 93;
  ram[1703]  = 195;
  ram[1704]  = 97;
  ram[1705]  = 14;
  ram[1706]  = 160;
  ram[1707]  = 209;
  ram[1708]  = 62;
  ram[1709]  = 53;
  ram[1710]  = 63;
  ram[1711]  = 61;
  ram[1712]  = 56;
  ram[1713]  = 52;
  ram[1714]  = 203;
  ram[1715]  = 164;
  ram[1716]  = 32;
  ram[1717]  = 57;
  ram[1718]  = 57;
  ram[1719]  = 61;
  ram[1720]  = 61;
  ram[1721]  = 67;
  ram[1722]  = 64;
  ram[1723]  = 68;
  ram[1724]  = 63;
  ram[1725]  = 64;
  ram[1726]  = 65;
  ram[1727]  = 65;
  ram[1728]  = 59;
  ram[1729]  = 66;
  ram[1730]  = 57;
  ram[1731]  = 62;
  ram[1732]  = 67;
  ram[1733]  = 61;
  ram[1734]  = 61;
  ram[1735]  = 58;
  ram[1736]  = 62;
  ram[1737]  = 52;
  ram[1738]  = 59;
  ram[1739]  = 32;
  ram[1740]  = 143;
  ram[1741]  = 207;
  ram[1742]  = 64;
  ram[1743]  = 13;
  ram[1744]  = 197;
  ram[1745]  = 203;
  ram[1746]  = 33;
  ram[1747]  = 58;
  ram[1748]  = 70;
  ram[1749]  = 55;
  ram[1750]  = 17;
  ram[1751]  = 74;
  ram[1752]  = 207;
  ram[1753]  = 121;
  ram[1754]  = 22;
  ram[1755]  = 128;
  ram[1756]  = 197;
  ram[1757]  = 75;
  ram[1758]  = 60;
  ram[1759]  = 64;
  ram[1760]  = 71;
  ram[1761]  = 58;
  ram[1762]  = 76;
  ram[1763]  = 186;
  ram[1764]  = 157;
  ram[1765]  = 23;
  ram[1766]  = 92;
  ram[1767]  = 200;
  ram[1768]  = 104;
  ram[1769]  = 43;
  ram[1770]  = 37;
  ram[1771]  = 0;
  ram[1772]  = 191;
  ram[1773]  = 224;
  ram[1774]  = 49;
  ram[1775]  = 54;
  ram[1776]  = 64;
  ram[1777]  = 43;
  ram[1778]  = 204;
  ram[1779]  = 167;
  ram[1780]  = 20;
  ram[1781]  = 60;
  ram[1782]  = 61;
  ram[1783]  = 58;
  ram[1784]  = 65;
  ram[1785]  = 62;
  ram[1786]  = 60;
  ram[1787]  = 66;
  ram[1788]  = 62;
  ram[1789]  = 65;
  ram[1790]  = 62;
  ram[1791]  = 64;
  ram[1792]  = 65;
  ram[1793]  = 60;
  ram[1794]  = 72;
  ram[1795]  = 62;
  ram[1796]  = 61;
  ram[1797]  = 74;
  ram[1798]  = 71;
  ram[1799]  = 80;
  ram[1800]  = 74;
  ram[1801]  = 72;
  ram[1802]  = 74;
  ram[1803]  = 64;
  ram[1804]  = 136;
  ram[1805]  = 201;
  ram[1806]  = 61;
  ram[1807]  = 17;
  ram[1808]  = 189;
  ram[1809]  = 197;
  ram[1810]  = 32;
  ram[1811]  = 59;
  ram[1812]  = 54;
  ram[1813]  = 67;
  ram[1814]  = 53;
  ram[1815]  = 93;
  ram[1816]  = 206;
  ram[1817]  = 112;
  ram[1818]  = 23;
  ram[1819]  = 129;
  ram[1820]  = 189;
  ram[1821]  = 78;
  ram[1822]  = 51;
  ram[1823]  = 67;
  ram[1824]  = 64;
  ram[1825]  = 67;
  ram[1826]  = 67;
  ram[1827]  = 190;
  ram[1828]  = 144;
  ram[1829]  = 29;
  ram[1830]  = 89;
  ram[1831]  = 205;
  ram[1832]  = 105;
  ram[1833]  = 47;
  ram[1834]  = 53;
  ram[1835]  = 36;
  ram[1836]  = 163;
  ram[1837]  = 187;
  ram[1838]  = 56;
  ram[1839]  = 84;
  ram[1840]  = 51;
  ram[1841]  = 40;
  ram[1842]  = 208;
  ram[1843]  = 151;
  ram[1844]  = 49;
  ram[1845]  = 66;
  ram[1846]  = 72;
  ram[1847]  = 66;
  ram[1848]  = 75;
  ram[1849]  = 79;
  ram[1850]  = 83;
  ram[1851]  = 63;
  ram[1852]  = 64;
  ram[1853]  = 61;
  ram[1854]  = 66;
  ram[1855]  = 67;
  ram[1856]  = 67;
  ram[1857]  = 66;
  ram[1858]  = 62;
  ram[1859]  = 65;
  ram[1860]  = 76;
  ram[1861]  = 212;
  ram[1862]  = 211;
  ram[1863]  = 209;
  ram[1864]  = 206;
  ram[1865]  = 211;
  ram[1866]  = 204;
  ram[1867]  = 221;
  ram[1868]  = 73;
  ram[1869]  = 19;
  ram[1870]  = 61;
  ram[1871]  = 23;
  ram[1872]  = 208;
  ram[1873]  = 202;
  ram[1874]  = 35;
  ram[1875]  = 62;
  ram[1876]  = 64;
  ram[1877]  = 60;
  ram[1878]  = 58;
  ram[1879]  = 104;
  ram[1880]  = 207;
  ram[1881]  = 130;
  ram[1882]  = 18;
  ram[1883]  = 142;
  ram[1884]  = 206;
  ram[1885]  = 85;
  ram[1886]  = 57;
  ram[1887]  = 69;
  ram[1888]  = 63;
  ram[1889]  = 67;
  ram[1890]  = 83;
  ram[1891]  = 200;
  ram[1892]  = 156;
  ram[1893]  = 23;
  ram[1894]  = 106;
  ram[1895]  = 214;
  ram[1896]  = 114;
  ram[1897]  = 48;
  ram[1898]  = 61;
  ram[1899]  = 60;
  ram[1900]  = 37;
  ram[1901]  = 0;
  ram[1902]  = 222;
  ram[1903]  = 228;
  ram[1904]  = 10;
  ram[1905]  = 50;
  ram[1906]  = 211;
  ram[1907]  = 186;
  ram[1908]  = 204;
  ram[1909]  = 205;
  ram[1910]  = 202;
  ram[1911]  = 206;
  ram[1912]  = 209;
  ram[1913]  = 209;
  ram[1914]  = 215;
  ram[1915]  = 95;
  ram[1916]  = 55;
  ram[1917]  = 61;
  ram[1918]  = 68;
  ram[1919]  = 63;
  ram[1920]  = 67;
  ram[1921]  = 69;
  ram[1922]  = 72;
  ram[1923]  = 62;
  ram[1924]  = 68;
  ram[1925]  = 161;
  ram[1926]  = 132;
  ram[1927]  = 155;
  ram[1928]  = 139;
  ram[1929]  = 156;
  ram[1930]  = 138;
  ram[1931]  = 166;
  ram[1932]  = 79;
  ram[1933]  = 55;
  ram[1934]  = 55;
  ram[1935]  = 46;
  ram[1936]  = 154;
  ram[1937]  = 163;
  ram[1938]  = 45;
  ram[1939]  = 56;
  ram[1940]  = 59;
  ram[1941]  = 68;
  ram[1942]  = 60;
  ram[1943]  = 89;
  ram[1944]  = 181;
  ram[1945]  = 93;
  ram[1946]  = 38;
  ram[1947]  = 114;
  ram[1948]  = 158;
  ram[1949]  = 72;
  ram[1950]  = 58;
  ram[1951]  = 63;
  ram[1952]  = 68;
  ram[1953]  = 58;
  ram[1954]  = 66;
  ram[1955]  = 162;
  ram[1956]  = 125;
  ram[1957]  = 44;
  ram[1958]  = 90;
  ram[1959]  = 175;
  ram[1960]  = 95;
  ram[1961]  = 53;
  ram[1962]  = 54;
  ram[1963]  = 62;
  ram[1964]  = 60;
  ram[1965]  = 40;
  ram[1966]  = 162;
  ram[1967]  = 179;
  ram[1968]  = 29;
  ram[1969]  = 49;
  ram[1970]  = 174;
  ram[1971]  = 132;
  ram[1972]  = 150;
  ram[1973]  = 136;
  ram[1974]  = 150;
  ram[1975]  = 136;
  ram[1976]  = 153;
  ram[1977]  = 136;
  ram[1978]  = 156;
  ram[1979]  = 81;
  ram[1980]  = 59;
  ram[1981]  = 63;
  ram[1982]  = 63;
  ram[1983]  = 67;
  ram[1984]  = 68;
  ram[1985]  = 69;
  ram[1986]  = 69;
  ram[1987]  = 70;
  ram[1988]  = 62;
  ram[1989]  = 43;
  ram[1990]  = 40;
  ram[1991]  = 36;
  ram[1992]  = 34;
  ram[1993]  = 34;
  ram[1994]  = 37;
  ram[1995]  = 39;
  ram[1996]  = 52;
  ram[1997]  = 64;
  ram[1998]  = 68;
  ram[1999]  = 61;
  ram[2000]  = 45;
  ram[2001]  = 38;
  ram[2002]  = 65;
  ram[2003]  = 63;
  ram[2004]  = 65;
  ram[2005]  = 65;
  ram[2006]  = 69;
  ram[2007]  = 54;
  ram[2008]  = 36;
  ram[2009]  = 56;
  ram[2010]  = 62;
  ram[2011]  = 40;
  ram[2012]  = 40;
  ram[2013]  = 56;
  ram[2014]  = 64;
  ram[2015]  = 67;
  ram[2016]  = 63;
  ram[2017]  = 62;
  ram[2018]  = 61;
  ram[2019]  = 35;
  ram[2020]  = 47;
  ram[2021]  = 63;
  ram[2022]  = 59;
  ram[2023]  = 45;
  ram[2024]  = 56;
  ram[2025]  = 64;
  ram[2026]  = 65;
  ram[2027]  = 65;
  ram[2028]  = 64;
  ram[2029]  = 64;
  ram[2030]  = 44;
  ram[2031]  = 40;
  ram[2032]  = 65;
  ram[2033]  = 58;
  ram[2034]  = 36;
  ram[2035]  = 43;
  ram[2036]  = 34;
  ram[2037]  = 30;
  ram[2038]  = 35;
  ram[2039]  = 36;
  ram[2040]  = 36;
  ram[2041]  = 39;
  ram[2042]  = 36;
  ram[2043]  = 46;
  ram[2044]  = 65;
  ram[2045]  = 62;
  ram[2046]  = 62;
  ram[2047]  = 64;
  ram[2048]  = 69;
  ram[2049]  = 69;
  ram[2050]  = 68;
  ram[2051]  = 67;
  ram[2052]  = 66;
  ram[2053]  = 66;
  ram[2054]  = 65;
  ram[2055]  = 65;
  ram[2056]  = 65;
  ram[2057]  = 67;
  ram[2058]  = 66;
  ram[2059]  = 65;
  ram[2060]  = 65;
  ram[2061]  = 65;
  ram[2062]  = 64;
  ram[2063]  = 63;
  ram[2064]  = 64;
  ram[2065]  = 65;
  ram[2066]  = 65;
  ram[2067]  = 65;
  ram[2068]  = 65;
  ram[2069]  = 66;
  ram[2070]  = 66;
  ram[2071]  = 66;
  ram[2072]  = 66;
  ram[2073]  = 66;
  ram[2074]  = 66;
  ram[2075]  = 65;
  ram[2076]  = 65;
  ram[2077]  = 65;
  ram[2078]  = 66;
  ram[2079]  = 67;
  ram[2080]  = 68;
  ram[2081]  = 68;
  ram[2082]  = 67;
  ram[2083]  = 68;
  ram[2084]  = 68;
  ram[2085]  = 66;
  ram[2086]  = 67;
  ram[2087]  = 67;
  ram[2088]  = 67;
  ram[2089]  = 67;
  ram[2090]  = 66;
  ram[2091]  = 66;
  ram[2092]  = 66;
  ram[2093]  = 66;
  ram[2094]  = 66;
  ram[2095]  = 66;
  ram[2096]  = 58;
  ram[2097]  = 61;
  ram[2098]  = 65;
  ram[2099]  = 66;
  ram[2100]  = 65;
  ram[2101]  = 64;
  ram[2102]  = 64;
  ram[2103]  = 65;
  ram[2104]  = 66;
  ram[2105]  = 66;
  ram[2106]  = 66;
  ram[2107]  = 66;
  ram[2108]  = 63;
  ram[2109]  = 62;
  ram[2110]  = 61;
  ram[2111]  = 61;
  ram[2112]  = 67;
  ram[2113]  = 67;
  ram[2114]  = 66;
  ram[2115]  = 66;
  ram[2116]  = 66;
  ram[2117]  = 66;
  ram[2118]  = 66;
  ram[2119]  = 66;
  ram[2120]  = 65;
  ram[2121]  = 66;
  ram[2122]  = 66;
  ram[2123]  = 63;
  ram[2124]  = 64;
  ram[2125]  = 64;
  ram[2126]  = 64;
  ram[2127]  = 64;
  ram[2128]  = 66;
  ram[2129]  = 67;
  ram[2130]  = 67;
  ram[2131]  = 68;
  ram[2132]  = 68;
  ram[2133]  = 68;
  ram[2134]  = 67;
  ram[2135]  = 67;
  ram[2136]  = 66;
  ram[2137]  = 66;
  ram[2138]  = 66;
  ram[2139]  = 66;
  ram[2140]  = 66;
  ram[2141]  = 66;
  ram[2142]  = 66;
  ram[2143]  = 66;
  ram[2144]  = 67;
  ram[2145]  = 66;
  ram[2146]  = 67;
  ram[2147]  = 66;
  ram[2148]  = 65;
  ram[2149]  = 64;
  ram[2150]  = 64;
  ram[2151]  = 65;
  ram[2152]  = 66;
  ram[2153]  = 66;
  ram[2154]  = 66;
  ram[2155]  = 67;
  ram[2156]  = 67;
  ram[2157]  = 67;
  ram[2158]  = 69;
  ram[2159]  = 67;
  ram[2160]  = 64;
  ram[2161]  = 65;
  ram[2162]  = 66;
  ram[2163]  = 66;
  ram[2164]  = 66;
  ram[2165]  = 65;
  ram[2166]  = 65;
  ram[2167]  = 65;
  ram[2168]  = 65;
  ram[2169]  = 65;
  ram[2170]  = 65;
  ram[2171]  = 65;
  ram[2172]  = 64;
  ram[2173]  = 61;
  ram[2174]  = 62;
  ram[2175]  = 60;
  ram[2176]  = 69;
  ram[2177]  = 69;
  ram[2178]  = 68;
  ram[2179]  = 68;
  ram[2180]  = 68;
  ram[2181]  = 68;
  ram[2182]  = 68;
  ram[2183]  = 66;
  ram[2184]  = 67;
  ram[2185]  = 67;
  ram[2186]  = 66;
  ram[2187]  = 63;
  ram[2188]  = 64;
  ram[2189]  = 64;
  ram[2190]  = 65;
  ram[2191]  = 66;
  ram[2192]  = 68;
  ram[2193]  = 71;
  ram[2194]  = 71;
  ram[2195]  = 71;
  ram[2196]  = 72;
  ram[2197]  = 72;
  ram[2198]  = 71;
  ram[2199]  = 71;
  ram[2200]  = 70;
  ram[2201]  = 70;
  ram[2202]  = 69;
  ram[2203]  = 69;
  ram[2204]  = 69;
  ram[2205]  = 69;
  ram[2206]  = 69;
  ram[2207]  = 69;
  ram[2208]  = 68;
  ram[2209]  = 67;
  ram[2210]  = 67;
  ram[2211]  = 65;
  ram[2212]  = 65;
  ram[2213]  = 64;
  ram[2214]  = 65;
  ram[2215]  = 66;
  ram[2216]  = 67;
  ram[2217]  = 67;
  ram[2218]  = 67;
  ram[2219]  = 69;
  ram[2220]  = 69;
  ram[2221]  = 69;
  ram[2222]  = 70;
  ram[2223]  = 69;
  ram[2224]  = 71;
  ram[2225]  = 69;
  ram[2226]  = 67;
  ram[2227]  = 65;
  ram[2228]  = 66;
  ram[2229]  = 66;
  ram[2230]  = 66;
  ram[2231]  = 65;
  ram[2232]  = 65;
  ram[2233]  = 65;
  ram[2234]  = 65;
  ram[2235]  = 65;
  ram[2236]  = 64;
  ram[2237]  = 62;
  ram[2238]  = 62;
  ram[2239]  = 61;
  ram[2240]  = 68;
  ram[2241]  = 68;
  ram[2242]  = 68;
  ram[2243]  = 68;
  ram[2244]  = 67;
  ram[2245]  = 67;
  ram[2246]  = 66;
  ram[2247]  = 66;
  ram[2248]  = 68;
  ram[2249]  = 65;
  ram[2250]  = 66;
  ram[2251]  = 63;
  ram[2252]  = 65;
  ram[2253]  = 64;
  ram[2254]  = 65;
  ram[2255]  = 67;
  ram[2256]  = 68;
  ram[2257]  = 68;
  ram[2258]  = 70;
  ram[2259]  = 69;
  ram[2260]  = 70;
  ram[2261]  = 69;
  ram[2262]  = 69;
  ram[2263]  = 69;
  ram[2264]  = 71;
  ram[2265]  = 69;
  ram[2266]  = 71;
  ram[2267]  = 69;
  ram[2268]  = 69;
  ram[2269]  = 68;
  ram[2270]  = 69;
  ram[2271]  = 69;
  ram[2272]  = 68;
  ram[2273]  = 66;
  ram[2274]  = 66;
  ram[2275]  = 66;
  ram[2276]  = 64;
  ram[2277]  = 63;
  ram[2278]  = 64;
  ram[2279]  = 66;
  ram[2280]  = 66;
  ram[2281]  = 66;
  ram[2282]  = 68;
  ram[2283]  = 68;
  ram[2284]  = 69;
  ram[2285]  = 68;
  ram[2286]  = 68;
  ram[2287]  = 67;
  ram[2288]  = 70;
  ram[2289]  = 67;
  ram[2290]  = 65;
  ram[2291]  = 65;
  ram[2292]  = 66;
  ram[2293]  = 65;
  ram[2294]  = 66;
  ram[2295]  = 64;
  ram[2296]  = 65;
  ram[2297]  = 64;
  ram[2298]  = 64;
  ram[2299]  = 63;
  ram[2300]  = 63;
  ram[2301]  = 61;
  ram[2302]  = 62;
  ram[2303]  = 60;
  ram[2304]  = 67;
  ram[2305]  = 67;
  ram[2306]  = 67;
  ram[2307]  = 67;
  ram[2308]  = 67;
  ram[2309]  = 66;
  ram[2310]  = 66;
  ram[2311]  = 65;
  ram[2312]  = 66;
  ram[2313]  = 65;
  ram[2314]  = 66;
  ram[2315]  = 65;
  ram[2316]  = 66;
  ram[2317]  = 64;
  ram[2318]  = 65;
  ram[2319]  = 66;
  ram[2320]  = 66;
  ram[2321]  = 66;
  ram[2322]  = 68;
  ram[2323]  = 66;
  ram[2324]  = 68;
  ram[2325]  = 66;
  ram[2326]  = 66;
  ram[2327]  = 66;
  ram[2328]  = 67;
  ram[2329]  = 65;
  ram[2330]  = 66;
  ram[2331]  = 65;
  ram[2332]  = 65;
  ram[2333]  = 65;
  ram[2334]  = 65;
  ram[2335]  = 65;
  ram[2336]  = 64;
  ram[2337]  = 63;
  ram[2338]  = 62;
  ram[2339]  = 62;
  ram[2340]  = 62;
  ram[2341]  = 62;
  ram[2342]  = 62;
  ram[2343]  = 64;
  ram[2344]  = 65;
  ram[2345]  = 65;
  ram[2346]  = 66;
  ram[2347]  = 66;
  ram[2348]  = 66;
  ram[2349]  = 66;
  ram[2350]  = 67;
  ram[2351]  = 65;
  ram[2352]  = 66;
  ram[2353]  = 65;
  ram[2354]  = 65;
  ram[2355]  = 65;
  ram[2356]  = 65;
  ram[2357]  = 64;
  ram[2358]  = 65;
  ram[2359]  = 64;
  ram[2360]  = 65;
  ram[2361]  = 64;
  ram[2362]  = 64;
  ram[2363]  = 62;
  ram[2364]  = 64;
  ram[2365]  = 61;
  ram[2366]  = 62;
  ram[2367]  = 59;
  ram[2368]  = 65;
  ram[2369]  = 65;
  ram[2370]  = 66;
  ram[2371]  = 66;
  ram[2372]  = 67;
  ram[2373]  = 66;
  ram[2374]  = 66;
  ram[2375]  = 65;
  ram[2376]  = 65;
  ram[2377]  = 65;
  ram[2378]  = 65;
  ram[2379]  = 66;
  ram[2380]  = 66;
  ram[2381]  = 65;
  ram[2382]  = 65;
  ram[2383]  = 65;
  ram[2384]  = 68;
  ram[2385]  = 68;
  ram[2386]  = 68;
  ram[2387]  = 68;
  ram[2388]  = 68;
  ram[2389]  = 66;
  ram[2390]  = 66;
  ram[2391]  = 66;
  ram[2392]  = 64;
  ram[2393]  = 63;
  ram[2394]  = 64;
  ram[2395]  = 63;
  ram[2396]  = 63;
  ram[2397]  = 61;
  ram[2398]  = 64;
  ram[2399]  = 64;
  ram[2400]  = 65;
  ram[2401]  = 64;
  ram[2402]  = 63;
  ram[2403]  = 64;
  ram[2404]  = 64;
  ram[2405]  = 63;
  ram[2406]  = 63;
  ram[2407]  = 64;
  ram[2408]  = 65;
  ram[2409]  = 65;
  ram[2410]  = 67;
  ram[2411]  = 68;
  ram[2412]  = 68;
  ram[2413]  = 68;
  ram[2414]  = 69;
  ram[2415]  = 68;
  ram[2416]  = 64;
  ram[2417]  = 65;
  ram[2418]  = 66;
  ram[2419]  = 66;
  ram[2420]  = 66;
  ram[2421]  = 65;
  ram[2422]  = 65;
  ram[2423]  = 65;
  ram[2424]  = 65;
  ram[2425]  = 65;
  ram[2426]  = 65;
  ram[2427]  = 64;
  ram[2428]  = 65;
  ram[2429]  = 63;
  ram[2430]  = 63;
  ram[2431]  = 62;
  ram[2432]  = 63;
  ram[2433]  = 64;
  ram[2434]  = 65;
  ram[2435]  = 65;
  ram[2436]  = 66;
  ram[2437]  = 65;
  ram[2438]  = 67;
  ram[2439]  = 66;
  ram[2440]  = 66;
  ram[2441]  = 66;
  ram[2442]  = 66;
  ram[2443]  = 67;
  ram[2444]  = 67;
  ram[2445]  = 66;
  ram[2446]  = 66;
  ram[2447]  = 67;
  ram[2448]  = 67;
  ram[2449]  = 67;
  ram[2450]  = 67;
  ram[2451]  = 67;
  ram[2452]  = 67;
  ram[2453]  = 66;
  ram[2454]  = 66;
  ram[2455]  = 66;
  ram[2456]  = 65;
  ram[2457]  = 63;
  ram[2458]  = 65;
  ram[2459]  = 63;
  ram[2460]  = 63;
  ram[2461]  = 62;
  ram[2462]  = 64;
  ram[2463]  = 64;
  ram[2464]  = 66;
  ram[2465]  = 65;
  ram[2466]  = 65;
  ram[2467]  = 66;
  ram[2468]  = 67;
  ram[2469]  = 66;
  ram[2470]  = 66;
  ram[2471]  = 66;
  ram[2472]  = 66;
  ram[2473]  = 67;
  ram[2474]  = 67;
  ram[2475]  = 68;
  ram[2476]  = 69;
  ram[2477]  = 69;
  ram[2478]  = 69;
  ram[2479]  = 68;
  ram[2480]  = 64;
  ram[2481]  = 63;
  ram[2482]  = 65;
  ram[2483]  = 65;
  ram[2484]  = 65;
  ram[2485]  = 64;
  ram[2486]  = 64;
  ram[2487]  = 64;
  ram[2488]  = 66;
  ram[2489]  = 66;
  ram[2490]  = 66;
  ram[2491]  = 64;
  ram[2492]  = 66;
  ram[2493]  = 63;
  ram[2494]  = 64;
  ram[2495]  = 62;
  ram[2496]  = 62;
  ram[2497]  = 62;
  ram[2498]  = 63;
  ram[2499]  = 63;
  ram[2500]  = 63;
  ram[2501]  = 62;
  ram[2502]  = 63;
  ram[2503]  = 62;
  ram[2504]  = 64;
  ram[2505]  = 63;
  ram[2506]  = 63;
  ram[2507]  = 64;
  ram[2508]  = 64;
  ram[2509]  = 64;
  ram[2510]  = 64;
  ram[2511]  = 66;
  ram[2512]  = 64;
  ram[2513]  = 65;
  ram[2514]  = 65;
  ram[2515]  = 63;
  ram[2516]  = 63;
  ram[2517]  = 63;
  ram[2518]  = 63;
  ram[2519]  = 63;
  ram[2520]  = 62;
  ram[2521]  = 62;
  ram[2522]  = 63;
  ram[2523]  = 61;
  ram[2524]  = 61;
  ram[2525]  = 61;
  ram[2526]  = 62;
  ram[2527]  = 62;
  ram[2528]  = 63;
  ram[2529]  = 62;
  ram[2530]  = 63;
  ram[2531]  = 64;
  ram[2532]  = 65;
  ram[2533]  = 64;
  ram[2534]  = 64;
  ram[2535]  = 64;
  ram[2536]  = 65;
  ram[2537]  = 65;
  ram[2538]  = 65;
  ram[2539]  = 65;
  ram[2540]  = 65;
  ram[2541]  = 64;
  ram[2542]  = 65;
  ram[2543]  = 64;
  ram[2544]  = 60;
  ram[2545]  = 59;
  ram[2546]  = 60;
  ram[2547]  = 61;
  ram[2548]  = 62;
  ram[2549]  = 62;
  ram[2550]  = 62;
  ram[2551]  = 62;
  ram[2552]  = 62;
  ram[2553]  = 63;
  ram[2554]  = 63;
  ram[2555]  = 63;
  ram[2556]  = 63;
  ram[2557]  = 62;
  ram[2558]  = 61;
  ram[2559]  = 61;
  ram[2560]  = 61;
  ram[2561]  = 61;
  ram[2562]  = 63;
  ram[2563]  = 62;
  ram[2564]  = 62;
  ram[2565]  = 62;
  ram[2566]  = 62;
  ram[2567]  = 62;
  ram[2568]  = 61;
  ram[2569]  = 62;
  ram[2570]  = 63;
  ram[2571]  = 62;
  ram[2572]  = 62;
  ram[2573]  = 62;
  ram[2574]  = 63;
  ram[2575]  = 64;
  ram[2576]  = 63;
  ram[2577]  = 48;
  ram[2578]  = 49;
  ram[2579]  = 46;
  ram[2580]  = 45;
  ram[2581]  = 44;
  ram[2582]  = 47;
  ram[2583]  = 44;
  ram[2584]  = 43;
  ram[2585]  = 43;
  ram[2586]  = 44;
  ram[2587]  = 41;
  ram[2588]  = 44;
  ram[2589]  = 42;
  ram[2590]  = 43;
  ram[2591]  = 44;
  ram[2592]  = 41;
  ram[2593]  = 38;
  ram[2594]  = 44;
  ram[2595]  = 40;
  ram[2596]  = 45;
  ram[2597]  = 44;
  ram[2598]  = 38;
  ram[2599]  = 45;
  ram[2600]  = 40;
  ram[2601]  = 41;
  ram[2602]  = 44;
  ram[2603]  = 40;
  ram[2604]  = 44;
  ram[2605]  = 47;
  ram[2606]  = 38;
  ram[2607]  = 58;
  ram[2608]  = 58;
  ram[2609]  = 59;
  ram[2610]  = 59;
  ram[2611]  = 58;
  ram[2612]  = 61;
  ram[2613]  = 61;
  ram[2614]  = 62;
  ram[2615]  = 61;
  ram[2616]  = 61;
  ram[2617]  = 62;
  ram[2618]  = 63;
  ram[2619]  = 63;
  ram[2620]  = 63;
  ram[2621]  = 62;
  ram[2622]  = 61;
  ram[2623]  = 60;
  ram[2624]  = 62;
  ram[2625]  = 62;
  ram[2626]  = 62;
  ram[2627]  = 62;
  ram[2628]  = 61;
  ram[2629]  = 61;
  ram[2630]  = 61;
  ram[2631]  = 61;
  ram[2632]  = 61;
  ram[2633]  = 62;
  ram[2634]  = 62;
  ram[2635]  = 62;
  ram[2636]  = 62;
  ram[2637]  = 62;
  ram[2638]  = 62;
  ram[2639]  = 62;
  ram[2640]  = 63;
  ram[2641]  = 149;
  ram[2642]  = 145;
  ram[2643]  = 146;
  ram[2644]  = 146;
  ram[2645]  = 139;
  ram[2646]  = 137;
  ram[2647]  = 142;
  ram[2648]  = 139;
  ram[2649]  = 142;
  ram[2650]  = 135;
  ram[2651]  = 141;
  ram[2652]  = 135;
  ram[2653]  = 143;
  ram[2654]  = 136;
  ram[2655]  = 139;
  ram[2656]  = 136;
  ram[2657]  = 139;
  ram[2658]  = 139;
  ram[2659]  = 134;
  ram[2660]  = 140;
  ram[2661]  = 130;
  ram[2662]  = 146;
  ram[2663]  = 131;
  ram[2664]  = 139;
  ram[2665]  = 136;
  ram[2666]  = 134;
  ram[2667]  = 135;
  ram[2668]  = 137;
  ram[2669]  = 127;
  ram[2670]  = 146;
  ram[2671]  = 55;
  ram[2672]  = 58;
  ram[2673]  = 60;
  ram[2674]  = 62;
  ram[2675]  = 60;
  ram[2676]  = 59;
  ram[2677]  = 60;
  ram[2678]  = 59;
  ram[2679]  = 59;
  ram[2680]  = 60;
  ram[2681]  = 61;
  ram[2682]  = 61;
  ram[2683]  = 61;
  ram[2684]  = 61;
  ram[2685]  = 61;
  ram[2686]  = 60;
  ram[2687]  = 60;
  ram[2688]  = 61;
  ram[2689]  = 61;
  ram[2690]  = 61;
  ram[2691]  = 60;
  ram[2692]  = 60;
  ram[2693]  = 60;
  ram[2694]  = 60;
  ram[2695]  = 60;
  ram[2696]  = 60;
  ram[2697]  = 61;
  ram[2698]  = 60;
  ram[2699]  = 61;
  ram[2700]  = 61;
  ram[2701]  = 61;
  ram[2702]  = 61;
  ram[2703]  = 59;
  ram[2704]  = 64;
  ram[2705]  = 215;
  ram[2706]  = 222;
  ram[2707]  = 213;
  ram[2708]  = 209;
  ram[2709]  = 213;
  ram[2710]  = 214;
  ram[2711]  = 211;
  ram[2712]  = 210;
  ram[2713]  = 211;
  ram[2714]  = 207;
  ram[2715]  = 210;
  ram[2716]  = 207;
  ram[2717]  = 211;
  ram[2718]  = 207;
  ram[2719]  = 207;
  ram[2720]  = 209;
  ram[2721]  = 205;
  ram[2722]  = 210;
  ram[2723]  = 208;
  ram[2724]  = 208;
  ram[2725]  = 208;
  ram[2726]  = 209;
  ram[2727]  = 213;
  ram[2728]  = 207;
  ram[2729]  = 203;
  ram[2730]  = 207;
  ram[2731]  = 209;
  ram[2732]  = 203;
  ram[2733]  = 191;
  ram[2734]  = 188;
  ram[2735]  = 58;
  ram[2736]  = 55;
  ram[2737]  = 58;
  ram[2738]  = 60;
  ram[2739]  = 60;
  ram[2740]  = 59;
  ram[2741]  = 59;
  ram[2742]  = 59;
  ram[2743]  = 60;
  ram[2744]  = 60;
  ram[2745]  = 61;
  ram[2746]  = 60;
  ram[2747]  = 60;
  ram[2748]  = 60;
  ram[2749]  = 60;
  ram[2750]  = 61;
  ram[2751]  = 61;
  ram[2752]  = 59;
  ram[2753]  = 59;
  ram[2754]  = 59;
  ram[2755]  = 59;
  ram[2756]  = 59;
  ram[2757]  = 58;
  ram[2758]  = 58;
  ram[2759]  = 58;
  ram[2760]  = 58;
  ram[2761]  = 58;
  ram[2762]  = 60;
  ram[2763]  = 58;
  ram[2764]  = 61;
  ram[2765]  = 59;
  ram[2766]  = 61;
  ram[2767]  = 58;
  ram[2768]  = 53;
  ram[2769]  = 87;
  ram[2770]  = 74;
  ram[2771]  = 78;
  ram[2772]  = 80;
  ram[2773]  = 73;
  ram[2774]  = 75;
  ram[2775]  = 76;
  ram[2776]  = 72;
  ram[2777]  = 76;
  ram[2778]  = 65;
  ram[2779]  = 80;
  ram[2780]  = 66;
  ram[2781]  = 78;
  ram[2782]  = 67;
  ram[2783]  = 70;
  ram[2784]  = 71;
  ram[2785]  = 79;
  ram[2786]  = 73;
  ram[2787]  = 68;
  ram[2788]  = 79;
  ram[2789]  = 70;
  ram[2790]  = 78;
  ram[2791]  = 69;
  ram[2792]  = 78;
  ram[2793]  = 67;
  ram[2794]  = 76;
  ram[2795]  = 62;
  ram[2796]  = 64;
  ram[2797]  = 169;
  ram[2798]  = 185;
  ram[2799]  = 52;
  ram[2800]  = 53;
  ram[2801]  = 57;
  ram[2802]  = 59;
  ram[2803]  = 58;
  ram[2804]  = 57;
  ram[2805]  = 58;
  ram[2806]  = 59;
  ram[2807]  = 60;
  ram[2808]  = 59;
  ram[2809]  = 59;
  ram[2810]  = 60;
  ram[2811]  = 58;
  ram[2812]  = 60;
  ram[2813]  = 58;
  ram[2814]  = 60;
  ram[2815]  = 59;
  ram[2816]  = 61;
  ram[2817]  = 61;
  ram[2818]  = 61;
  ram[2819]  = 60;
  ram[2820]  = 60;
  ram[2821]  = 60;
  ram[2822]  = 60;
  ram[2823]  = 60;
  ram[2824]  = 59;
  ram[2825]  = 60;
  ram[2826]  = 61;
  ram[2827]  = 60;
  ram[2828]  = 61;
  ram[2829]  = 59;
  ram[2830]  = 60;
  ram[2831]  = 61;
  ram[2832]  = 60;
  ram[2833]  = 46;
  ram[2834]  = 52;
  ram[2835]  = 49;
  ram[2836]  = 47;
  ram[2837]  = 42;
  ram[2838]  = 49;
  ram[2839]  = 46;
  ram[2840]  = 47;
  ram[2841]  = 45;
  ram[2842]  = 48;
  ram[2843]  = 46;
  ram[2844]  = 46;
  ram[2845]  = 43;
  ram[2846]  = 47;
  ram[2847]  = 44;
  ram[2848]  = 54;
  ram[2849]  = 46;
  ram[2850]  = 50;
  ram[2851]  = 51;
  ram[2852]  = 49;
  ram[2853]  = 51;
  ram[2854]  = 54;
  ram[2855]  = 45;
  ram[2856]  = 48;
  ram[2857]  = 48;
  ram[2858]  = 41;
  ram[2859]  = 39;
  ram[2860]  = 26;
  ram[2861]  = 183;
  ram[2862]  = 188;
  ram[2863]  = 55;
  ram[2864]  = 56;
  ram[2865]  = 59;
  ram[2866]  = 61;
  ram[2867]  = 60;
  ram[2868]  = 59;
  ram[2869]  = 59;
  ram[2870]  = 60;
  ram[2871]  = 60;
  ram[2872]  = 59;
  ram[2873]  = 59;
  ram[2874]  = 61;
  ram[2875]  = 60;
  ram[2876]  = 61;
  ram[2877]  = 59;
  ram[2878]  = 59;
  ram[2879]  = 58;
  ram[2880]  = 65;
  ram[2881]  = 63;
  ram[2882]  = 64;
  ram[2883]  = 62;
  ram[2884]  = 64;
  ram[2885]  = 61;
  ram[2886]  = 63;
  ram[2887]  = 61;
  ram[2888]  = 64;
  ram[2889]  = 63;
  ram[2890]  = 65;
  ram[2891]  = 62;
  ram[2892]  = 63;
  ram[2893]  = 60;
  ram[2894]  = 62;
  ram[2895]  = 62;
  ram[2896]  = 65;
  ram[2897]  = 60;
  ram[2898]  = 64;
  ram[2899]  = 60;
  ram[2900]  = 63;
  ram[2901]  = 61;
  ram[2902]  = 62;
  ram[2903]  = 61;
  ram[2904]  = 61;
  ram[2905]  = 61;
  ram[2906]  = 60;
  ram[2907]  = 63;
  ram[2908]  = 57;
  ram[2909]  = 64;
  ram[2910]  = 64;
  ram[2911]  = 61;
  ram[2912]  = 56;
  ram[2913]  = 62;
  ram[2914]  = 64;
  ram[2915]  = 64;
  ram[2916]  = 66;
  ram[2917]  = 60;
  ram[2918]  = 61;
  ram[2919]  = 61;
  ram[2920]  = 62;
  ram[2921]  = 57;
  ram[2922]  = 55;
  ram[2923]  = 41;
  ram[2924]  = 37;
  ram[2925]  = 179;
  ram[2926]  = 187;
  ram[2927]  = 54;
  ram[2928]  = 57;
  ram[2929]  = 60;
  ram[2930]  = 64;
  ram[2931]  = 61;
  ram[2932]  = 63;
  ram[2933]  = 61;
  ram[2934]  = 64;
  ram[2935]  = 62;
  ram[2936]  = 63;
  ram[2937]  = 61;
  ram[2938]  = 64;
  ram[2939]  = 62;
  ram[2940]  = 64;
  ram[2941]  = 61;
  ram[2942]  = 62;
  ram[2943]  = 60;
  ram[2944]  = 65;
  ram[2945]  = 64;
  ram[2946]  = 65;
  ram[2947]  = 63;
  ram[2948]  = 64;
  ram[2949]  = 63;
  ram[2950]  = 63;
  ram[2951]  = 62;
  ram[2952]  = 65;
  ram[2953]  = 63;
  ram[2954]  = 64;
  ram[2955]  = 62;
  ram[2956]  = 63;
  ram[2957]  = 61;
  ram[2958]  = 62;
  ram[2959]  = 62;
  ram[2960]  = 61;
  ram[2961]  = 69;
  ram[2962]  = 65;
  ram[2963]  = 63;
  ram[2964]  = 65;
  ram[2965]  = 64;
  ram[2966]  = 60;
  ram[2967]  = 60;
  ram[2968]  = 63;
  ram[2969]  = 59;
  ram[2970]  = 64;
  ram[2971]  = 59;
  ram[2972]  = 64;
  ram[2973]  = 64;
  ram[2974]  = 66;
  ram[2975]  = 52;
  ram[2976]  = 76;
  ram[2977]  = 71;
  ram[2978]  = 57;
  ram[2979]  = 63;
  ram[2980]  = 63;
  ram[2981]  = 64;
  ram[2982]  = 59;
  ram[2983]  = 61;
  ram[2984]  = 67;
  ram[2985]  = 59;
  ram[2986]  = 54;
  ram[2987]  = 55;
  ram[2988]  = 38;
  ram[2989]  = 182;
  ram[2990]  = 192;
  ram[2991]  = 47;
  ram[2992]  = 56;
  ram[2993]  = 60;
  ram[2994]  = 63;
  ram[2995]  = 62;
  ram[2996]  = 64;
  ram[2997]  = 63;
  ram[2998]  = 65;
  ram[2999]  = 63;
  ram[3000]  = 64;
  ram[3001]  = 63;
  ram[3002]  = 64;
  ram[3003]  = 63;
  ram[3004]  = 64;
  ram[3005]  = 63;
  ram[3006]  = 63;
  ram[3007]  = 62;
  ram[3008]  = 65;
  ram[3009]  = 64;
  ram[3010]  = 64;
  ram[3011]  = 64;
  ram[3012]  = 63;
  ram[3013]  = 63;
  ram[3014]  = 63;
  ram[3015]  = 63;
  ram[3016]  = 63;
  ram[3017]  = 62;
  ram[3018]  = 62;
  ram[3019]  = 62;
  ram[3020]  = 62;
  ram[3021]  = 63;
  ram[3022]  = 63;
  ram[3023]  = 62;
  ram[3024]  = 65;
  ram[3025]  = 63;
  ram[3026]  = 62;
  ram[3027]  = 66;
  ram[3028]  = 63;
  ram[3029]  = 63;
  ram[3030]  = 63;
  ram[3031]  = 64;
  ram[3032]  = 65;
  ram[3033]  = 62;
  ram[3034]  = 63;
  ram[3035]  = 63;
  ram[3036]  = 62;
  ram[3037]  = 65;
  ram[3038]  = 57;
  ram[3039]  = 37;
  ram[3040]  = 251;
  ram[3041]  = 247;
  ram[3042]  = 33;
  ram[3043]  = 64;
  ram[3044]  = 65;
  ram[3045]  = 60;
  ram[3046]  = 49;
  ram[3047]  = 147;
  ram[3048]  = 219;
  ram[3049]  = 194;
  ram[3050]  = 200;
  ram[3051]  = 195;
  ram[3052]  = 193;
  ram[3053]  = 183;
  ram[3054]  = 193;
  ram[3055]  = 57;
  ram[3056]  = 59;
  ram[3057]  = 62;
  ram[3058]  = 63;
  ram[3059]  = 63;
  ram[3060]  = 63;
  ram[3061]  = 63;
  ram[3062]  = 62;
  ram[3063]  = 61;
  ram[3064]  = 62;
  ram[3065]  = 62;
  ram[3066]  = 62;
  ram[3067]  = 62;
  ram[3068]  = 62;
  ram[3069]  = 62;
  ram[3070]  = 63;
  ram[3071]  = 63;
  ram[3072]  = 66;
  ram[3073]  = 66;
  ram[3074]  = 67;
  ram[3075]  = 67;
  ram[3076]  = 67;
  ram[3077]  = 67;
  ram[3078]  = 66;
  ram[3079]  = 66;
  ram[3080]  = 67;
  ram[3081]  = 67;
  ram[3082]  = 67;
  ram[3083]  = 67;
  ram[3084]  = 67;
  ram[3085]  = 67;
  ram[3086]  = 67;
  ram[3087]  = 67;
  ram[3088]  = 68;
  ram[3089]  = 67;
  ram[3090]  = 66;
  ram[3091]  = 67;
  ram[3092]  = 68;
  ram[3093]  = 69;
  ram[3094]  = 68;
  ram[3095]  = 66;
  ram[3096]  = 69;
  ram[3097]  = 68;
  ram[3098]  = 68;
  ram[3099]  = 69;
  ram[3100]  = 66;
  ram[3101]  = 71;
  ram[3102]  = 68;
  ram[3103]  = 42;
  ram[3104]  = 234;
  ram[3105]  = 218;
  ram[3106]  = 35;
  ram[3107]  = 63;
  ram[3108]  = 63;
  ram[3109]  = 63;
  ram[3110]  = 48;
  ram[3111]  = 125;
  ram[3112]  = 196;
  ram[3113]  = 187;
  ram[3114]  = 184;
  ram[3115]  = 179;
  ram[3116]  = 180;
  ram[3117]  = 179;
  ram[3118]  = 174;
  ram[3119]  = 62;
  ram[3120]  = 61;
  ram[3121]  = 63;
  ram[3122]  = 63;
  ram[3123]  = 64;
  ram[3124]  = 64;
  ram[3125]  = 65;
  ram[3126]  = 67;
  ram[3127]  = 67;
  ram[3128]  = 67;
  ram[3129]  = 67;
  ram[3130]  = 67;
  ram[3131]  = 66;
  ram[3132]  = 66;
  ram[3133]  = 66;
  ram[3134]  = 68;
  ram[3135]  = 67;
  ram[3136]  = 69;
  ram[3137]  = 69;
  ram[3138]  = 69;
  ram[3139]  = 70;
  ram[3140]  = 70;
  ram[3141]  = 69;
  ram[3142]  = 69;
  ram[3143]  = 69;
  ram[3144]  = 68;
  ram[3145]  = 68;
  ram[3146]  = 68;
  ram[3147]  = 68;
  ram[3148]  = 68;
  ram[3149]  = 68;
  ram[3150]  = 69;
  ram[3151]  = 69;
  ram[3152]  = 69;
  ram[3153]  = 68;
  ram[3154]  = 68;
  ram[3155]  = 68;
  ram[3156]  = 70;
  ram[3157]  = 70;
  ram[3158]  = 69;
  ram[3159]  = 68;
  ram[3160]  = 68;
  ram[3161]  = 68;
  ram[3162]  = 69;
  ram[3163]  = 71;
  ram[3164]  = 67;
  ram[3165]  = 69;
  ram[3166]  = 72;
  ram[3167]  = 59;
  ram[3168]  = 63;
  ram[3169]  = 56;
  ram[3170]  = 66;
  ram[3171]  = 66;
  ram[3172]  = 64;
  ram[3173]  = 67;
  ram[3174]  = 61;
  ram[3175]  = 56;
  ram[3176]  = 45;
  ram[3177]  = 45;
  ram[3178]  = 49;
  ram[3179]  = 44;
  ram[3180]  = 51;
  ram[3181]  = 44;
  ram[3182]  = 53;
  ram[3183]  = 59;
  ram[3184]  = 65;
  ram[3185]  = 65;
  ram[3186]  = 66;
  ram[3187]  = 66;
  ram[3188]  = 66;
  ram[3189]  = 67;
  ram[3190]  = 69;
  ram[3191]  = 69;
  ram[3192]  = 68;
  ram[3193]  = 69;
  ram[3194]  = 69;
  ram[3195]  = 68;
  ram[3196]  = 68;
  ram[3197]  = 68;
  ram[3198]  = 69;
  ram[3199]  = 68;
  ram[3200]  = 70;
  ram[3201]  = 70;
  ram[3202]  = 70;
  ram[3203]  = 70;
  ram[3204]  = 70;
  ram[3205]  = 69;
  ram[3206]  = 69;
  ram[3207]  = 69;
  ram[3208]  = 69;
  ram[3209]  = 68;
  ram[3210]  = 68;
  ram[3211]  = 68;
  ram[3212]  = 69;
  ram[3213]  = 69;
  ram[3214]  = 69;
  ram[3215]  = 69;
  ram[3216]  = 69;
  ram[3217]  = 68;
  ram[3218]  = 68;
  ram[3219]  = 68;
  ram[3220]  = 69;
  ram[3221]  = 70;
  ram[3222]  = 69;
  ram[3223]  = 68;
  ram[3224]  = 67;
  ram[3225]  = 67;
  ram[3226]  = 68;
  ram[3227]  = 70;
  ram[3228]  = 68;
  ram[3229]  = 67;
  ram[3230]  = 72;
  ram[3231]  = 70;
  ram[3232]  = 59;
  ram[3233]  = 65;
  ram[3234]  = 65;
  ram[3235]  = 66;
  ram[3236]  = 69;
  ram[3237]  = 63;
  ram[3238]  = 63;
  ram[3239]  = 57;
  ram[3240]  = 66;
  ram[3241]  = 56;
  ram[3242]  = 61;
  ram[3243]  = 56;
  ram[3244]  = 55;
  ram[3245]  = 63;
  ram[3246]  = 61;
  ram[3247]  = 67;
  ram[3248]  = 65;
  ram[3249]  = 67;
  ram[3250]  = 67;
  ram[3251]  = 67;
  ram[3252]  = 68;
  ram[3253]  = 68;
  ram[3254]  = 69;
  ram[3255]  = 69;
  ram[3256]  = 69;
  ram[3257]  = 70;
  ram[3258]  = 70;
  ram[3259]  = 69;
  ram[3260]  = 69;
  ram[3261]  = 69;
  ram[3262]  = 69;
  ram[3263]  = 68;
  ram[3264]  = 70;
  ram[3265]  = 70;
  ram[3266]  = 70;
  ram[3267]  = 70;
  ram[3268]  = 69;
  ram[3269]  = 69;
  ram[3270]  = 69;
  ram[3271]  = 69;
  ram[3272]  = 69;
  ram[3273]  = 69;
  ram[3274]  = 69;
  ram[3275]  = 69;
  ram[3276]  = 70;
  ram[3277]  = 70;
  ram[3278]  = 70;
  ram[3279]  = 70;
  ram[3280]  = 70;
  ram[3281]  = 69;
  ram[3282]  = 69;
  ram[3283]  = 69;
  ram[3284]  = 70;
  ram[3285]  = 70;
  ram[3286]  = 69;
  ram[3287]  = 68;
  ram[3288]  = 69;
  ram[3289]  = 69;
  ram[3290]  = 67;
  ram[3291]  = 69;
  ram[3292]  = 70;
  ram[3293]  = 69;
  ram[3294]  = 69;
  ram[3295]  = 69;
  ram[3296]  = 71;
  ram[3297]  = 69;
  ram[3298]  = 67;
  ram[3299]  = 73;
  ram[3300]  = 66;
  ram[3301]  = 66;
  ram[3302]  = 70;
  ram[3303]  = 67;
  ram[3304]  = 61;
  ram[3305]  = 66;
  ram[3306]  = 66;
  ram[3307]  = 68;
  ram[3308]  = 66;
  ram[3309]  = 68;
  ram[3310]  = 68;
  ram[3311]  = 70;
  ram[3312]  = 67;
  ram[3313]  = 67;
  ram[3314]  = 68;
  ram[3315]  = 68;
  ram[3316]  = 69;
  ram[3317]  = 69;
  ram[3318]  = 70;
  ram[3319]  = 71;
  ram[3320]  = 70;
  ram[3321]  = 71;
  ram[3322]  = 70;
  ram[3323]  = 70;
  ram[3324]  = 69;
  ram[3325]  = 69;
  ram[3326]  = 69;
  ram[3327]  = 68;
  ram[3328]  = 71;
  ram[3329]  = 71;
  ram[3330]  = 71;
  ram[3331]  = 71;
  ram[3332]  = 71;
  ram[3333]  = 71;
  ram[3334]  = 71;
  ram[3335]  = 71;
  ram[3336]  = 71;
  ram[3337]  = 71;
  ram[3338]  = 71;
  ram[3339]  = 71;
  ram[3340]  = 71;
  ram[3341]  = 71;
  ram[3342]  = 71;
  ram[3343]  = 71;
  ram[3344]  = 72;
  ram[3345]  = 72;
  ram[3346]  = 71;
  ram[3347]  = 72;
  ram[3348]  = 72;
  ram[3349]  = 72;
  ram[3350]  = 72;
  ram[3351]  = 71;
  ram[3352]  = 71;
  ram[3353]  = 73;
  ram[3354]  = 71;
  ram[3355]  = 70;
  ram[3356]  = 72;
  ram[3357]  = 72;
  ram[3358]  = 70;
  ram[3359]  = 70;
  ram[3360]  = 70;
  ram[3361]  = 71;
  ram[3362]  = 75;
  ram[3363]  = 69;
  ram[3364]  = 69;
  ram[3365]  = 73;
  ram[3366]  = 66;
  ram[3367]  = 71;
  ram[3368]  = 71;
  ram[3369]  = 67;
  ram[3370]  = 65;
  ram[3371]  = 72;
  ram[3372]  = 71;
  ram[3373]  = 66;
  ram[3374]  = 73;
  ram[3375]  = 69;
  ram[3376]  = 70;
  ram[3377]  = 70;
  ram[3378]  = 71;
  ram[3379]  = 71;
  ram[3380]  = 72;
  ram[3381]  = 71;
  ram[3382]  = 72;
  ram[3383]  = 72;
  ram[3384]  = 71;
  ram[3385]  = 71;
  ram[3386]  = 71;
  ram[3387]  = 70;
  ram[3388]  = 70;
  ram[3389]  = 70;
  ram[3390]  = 69;
  ram[3391]  = 68;
  ram[3392]  = 71;
  ram[3393]  = 71;
  ram[3394]  = 71;
  ram[3395]  = 71;
  ram[3396]  = 71;
  ram[3397]  = 72;
  ram[3398]  = 72;
  ram[3399]  = 72;
  ram[3400]  = 73;
  ram[3401]  = 73;
  ram[3402]  = 73;
  ram[3403]  = 73;
  ram[3404]  = 73;
  ram[3405]  = 73;
  ram[3406]  = 73;
  ram[3407]  = 72;
  ram[3408]  = 72;
  ram[3409]  = 72;
  ram[3410]  = 71;
  ram[3411]  = 72;
  ram[3412]  = 72;
  ram[3413]  = 72;
  ram[3414]  = 71;
  ram[3415]  = 71;
  ram[3416]  = 69;
  ram[3417]  = 72;
  ram[3418]  = 74;
  ram[3419]  = 70;
  ram[3420]  = 70;
  ram[3421]  = 72;
  ram[3422]  = 71;
  ram[3423]  = 74;
  ram[3424]  = 79;
  ram[3425]  = 74;
  ram[3426]  = 68;
  ram[3427]  = 80;
  ram[3428]  = 69;
  ram[3429]  = 72;
  ram[3430]  = 74;
  ram[3431]  = 70;
  ram[3432]  = 67;
  ram[3433]  = 75;
  ram[3434]  = 74;
  ram[3435]  = 68;
  ram[3436]  = 76;
  ram[3437]  = 70;
  ram[3438]  = 68;
  ram[3439]  = 77;
  ram[3440]  = 74;
  ram[3441]  = 73;
  ram[3442]  = 73;
  ram[3443]  = 72;
  ram[3444]  = 72;
  ram[3445]  = 72;
  ram[3446]  = 72;
  ram[3447]  = 72;
  ram[3448]  = 72;
  ram[3449]  = 73;
  ram[3450]  = 73;
  ram[3451]  = 72;
  ram[3452]  = 71;
  ram[3453]  = 71;
  ram[3454]  = 70;
  ram[3455]  = 69;
  ram[3456]  = 72;
  ram[3457]  = 72;
  ram[3458]  = 72;
  ram[3459]  = 72;
  ram[3460]  = 73;
  ram[3461]  = 73;
  ram[3462]  = 74;
  ram[3463]  = 74;
  ram[3464]  = 75;
  ram[3465]  = 75;
  ram[3466]  = 75;
  ram[3467]  = 75;
  ram[3468]  = 75;
  ram[3469]  = 74;
  ram[3470]  = 74;
  ram[3471]  = 73;
  ram[3472]  = 72;
  ram[3473]  = 72;
  ram[3474]  = 71;
  ram[3475]  = 71;
  ram[3476]  = 72;
  ram[3477]  = 71;
  ram[3478]  = 71;
  ram[3479]  = 70;
  ram[3480]  = 70;
  ram[3481]  = 70;
  ram[3482]  = 74;
  ram[3483]  = 72;
  ram[3484]  = 70;
  ram[3485]  = 73;
  ram[3486]  = 72;
  ram[3487]  = 75;
  ram[3488]  = 73;
  ram[3489]  = 72;
  ram[3490]  = 78;
  ram[3491]  = 74;
  ram[3492]  = 69;
  ram[3493]  = 72;
  ram[3494]  = 77;
  ram[3495]  = 71;
  ram[3496]  = 82;
  ram[3497]  = 69;
  ram[3498]  = 73;
  ram[3499]  = 76;
  ram[3500]  = 73;
  ram[3501]  = 73;
  ram[3502]  = 76;
  ram[3503]  = 75;
  ram[3504]  = 76;
  ram[3505]  = 75;
  ram[3506]  = 75;
  ram[3507]  = 75;
  ram[3508]  = 74;
  ram[3509]  = 74;
  ram[3510]  = 72;
  ram[3511]  = 72;
  ram[3512]  = 74;
  ram[3513]  = 75;
  ram[3514]  = 75;
  ram[3515]  = 74;
  ram[3516]  = 73;
  ram[3517]  = 73;
  ram[3518]  = 72;
  ram[3519]  = 71;
  ram[3520]  = 74;
  ram[3521]  = 73;
  ram[3522]  = 73;
  ram[3523]  = 74;
  ram[3524]  = 74;
  ram[3525]  = 75;
  ram[3526]  = 75;
  ram[3527]  = 76;
  ram[3528]  = 75;
  ram[3529]  = 75;
  ram[3530]  = 75;
  ram[3531]  = 75;
  ram[3532]  = 75;
  ram[3533]  = 74;
  ram[3534]  = 73;
  ram[3535]  = 73;
  ram[3536]  = 74;
  ram[3537]  = 73;
  ram[3538]  = 73;
  ram[3539]  = 73;
  ram[3540]  = 73;
  ram[3541]  = 73;
  ram[3542]  = 72;
  ram[3543]  = 72;
  ram[3544]  = 74;
  ram[3545]  = 70;
  ram[3546]  = 75;
  ram[3547]  = 75;
  ram[3548]  = 75;
  ram[3549]  = 76;
  ram[3550]  = 73;
  ram[3551]  = 73;
  ram[3552]  = 73;
  ram[3553]  = 78;
  ram[3554]  = 69;
  ram[3555]  = 75;
  ram[3556]  = 75;
  ram[3557]  = 73;
  ram[3558]  = 71;
  ram[3559]  = 73;
  ram[3560]  = 72;
  ram[3561]  = 78;
  ram[3562]  = 76;
  ram[3563]  = 74;
  ram[3564]  = 75;
  ram[3565]  = 78;
  ram[3566]  = 79;
  ram[3567]  = 75;
  ram[3568]  = 76;
  ram[3569]  = 76;
  ram[3570]  = 76;
  ram[3571]  = 76;
  ram[3572]  = 76;
  ram[3573]  = 76;
  ram[3574]  = 74;
  ram[3575]  = 75;
  ram[3576]  = 74;
  ram[3577]  = 75;
  ram[3578]  = 76;
  ram[3579]  = 75;
  ram[3580]  = 74;
  ram[3581]  = 74;
  ram[3582]  = 73;
  ram[3583]  = 71;
  ram[3584]  = 75;
  ram[3585]  = 75;
  ram[3586]  = 75;
  ram[3587]  = 74;
  ram[3588]  = 74;
  ram[3589]  = 74;
  ram[3590]  = 74;
  ram[3591]  = 73;
  ram[3592]  = 73;
  ram[3593]  = 73;
  ram[3594]  = 73;
  ram[3595]  = 73;
  ram[3596]  = 73;
  ram[3597]  = 73;
  ram[3598]  = 73;
  ram[3599]  = 73;
  ram[3600]  = 72;
  ram[3601]  = 72;
  ram[3602]  = 72;
  ram[3603]  = 73;
  ram[3604]  = 73;
  ram[3605]  = 73;
  ram[3606]  = 73;
  ram[3607]  = 73;
  ram[3608]  = 73;
  ram[3609]  = 73;
  ram[3610]  = 73;
  ram[3611]  = 73;
  ram[3612]  = 73;
  ram[3613]  = 73;
  ram[3614]  = 73;
  ram[3615]  = 73;
  ram[3616]  = 74;
  ram[3617]  = 73;
  ram[3618]  = 72;
  ram[3619]  = 72;
  ram[3620]  = 72;
  ram[3621]  = 72;
  ram[3622]  = 72;
  ram[3623]  = 72;
  ram[3624]  = 73;
  ram[3625]  = 73;
  ram[3626]  = 73;
  ram[3627]  = 73;
  ram[3628]  = 76;
  ram[3629]  = 76;
  ram[3630]  = 76;
  ram[3631]  = 76;
  ram[3632]  = 77;
  ram[3633]  = 77;
  ram[3634]  = 77;
  ram[3635]  = 77;
  ram[3636]  = 76;
  ram[3637]  = 76;
  ram[3638]  = 76;
  ram[3639]  = 76;
  ram[3640]  = 75;
  ram[3641]  = 75;
  ram[3642]  = 75;
  ram[3643]  = 75;
  ram[3644]  = 74;
  ram[3645]  = 73;
  ram[3646]  = 73;
  ram[3647]  = 72;
  ram[3648]  = 74;
  ram[3649]  = 75;
  ram[3650]  = 75;
  ram[3651]  = 74;
  ram[3652]  = 74;
  ram[3653]  = 75;
  ram[3654]  = 75;
  ram[3655]  = 74;
  ram[3656]  = 76;
  ram[3657]  = 76;
  ram[3658]  = 76;
  ram[3659]  = 76;
  ram[3660]  = 76;
  ram[3661]  = 76;
  ram[3662]  = 76;
  ram[3663]  = 76;
  ram[3664]  = 76;
  ram[3665]  = 76;
  ram[3666]  = 76;
  ram[3667]  = 76;
  ram[3668]  = 76;
  ram[3669]  = 76;
  ram[3670]  = 76;
  ram[3671]  = 76;
  ram[3672]  = 75;
  ram[3673]  = 75;
  ram[3674]  = 75;
  ram[3675]  = 75;
  ram[3676]  = 75;
  ram[3677]  = 75;
  ram[3678]  = 75;
  ram[3679]  = 75;
  ram[3680]  = 74;
  ram[3681]  = 74;
  ram[3682]  = 74;
  ram[3683]  = 74;
  ram[3684]  = 74;
  ram[3685]  = 74;
  ram[3686]  = 73;
  ram[3687]  = 73;
  ram[3688]  = 75;
  ram[3689]  = 75;
  ram[3690]  = 75;
  ram[3691]  = 75;
  ram[3692]  = 77;
  ram[3693]  = 77;
  ram[3694]  = 78;
  ram[3695]  = 78;
  ram[3696]  = 78;
  ram[3697]  = 78;
  ram[3698]  = 78;
  ram[3699]  = 78;
  ram[3700]  = 78;
  ram[3701]  = 78;
  ram[3702]  = 78;
  ram[3703]  = 78;
  ram[3704]  = 75;
  ram[3705]  = 75;
  ram[3706]  = 75;
  ram[3707]  = 75;
  ram[3708]  = 74;
  ram[3709]  = 73;
  ram[3710]  = 73;
  ram[3711]  = 72;
  ram[3712]  = 75;
  ram[3713]  = 75;
  ram[3714]  = 75;
  ram[3715]  = 74;
  ram[3716]  = 75;
  ram[3717]  = 76;
  ram[3718]  = 76;
  ram[3719]  = 76;
  ram[3720]  = 76;
  ram[3721]  = 76;
  ram[3722]  = 76;
  ram[3723]  = 76;
  ram[3724]  = 75;
  ram[3725]  = 75;
  ram[3726]  = 75;
  ram[3727]  = 75;
  ram[3728]  = 75;
  ram[3729]  = 75;
  ram[3730]  = 75;
  ram[3731]  = 75;
  ram[3732]  = 75;
  ram[3733]  = 75;
  ram[3734]  = 75;
  ram[3735]  = 75;
  ram[3736]  = 75;
  ram[3737]  = 75;
  ram[3738]  = 75;
  ram[3739]  = 75;
  ram[3740]  = 75;
  ram[3741]  = 75;
  ram[3742]  = 75;
  ram[3743]  = 75;
  ram[3744]  = 74;
  ram[3745]  = 74;
  ram[3746]  = 74;
  ram[3747]  = 74;
  ram[3748]  = 74;
  ram[3749]  = 73;
  ram[3750]  = 73;
  ram[3751]  = 73;
  ram[3752]  = 74;
  ram[3753]  = 74;
  ram[3754]  = 74;
  ram[3755]  = 74;
  ram[3756]  = 75;
  ram[3757]  = 75;
  ram[3758]  = 75;
  ram[3759]  = 76;
  ram[3760]  = 77;
  ram[3761]  = 77;
  ram[3762]  = 77;
  ram[3763]  = 77;
  ram[3764]  = 75;
  ram[3765]  = 75;
  ram[3766]  = 75;
  ram[3767]  = 75;
  ram[3768]  = 75;
  ram[3769]  = 75;
  ram[3770]  = 75;
  ram[3771]  = 75;
  ram[3772]  = 74;
  ram[3773]  = 73;
  ram[3774]  = 73;
  ram[3775]  = 72;
  ram[3776]  = 76;
  ram[3777]  = 76;
  ram[3778]  = 76;
  ram[3779]  = 75;
  ram[3780]  = 75;
  ram[3781]  = 76;
  ram[3782]  = 76;
  ram[3783]  = 76;
  ram[3784]  = 77;
  ram[3785]  = 76;
  ram[3786]  = 76;
  ram[3787]  = 76;
  ram[3788]  = 76;
  ram[3789]  = 76;
  ram[3790]  = 76;
  ram[3791]  = 76;
  ram[3792]  = 76;
  ram[3793]  = 76;
  ram[3794]  = 76;
  ram[3795]  = 76;
  ram[3796]  = 76;
  ram[3797]  = 76;
  ram[3798]  = 76;
  ram[3799]  = 76;
  ram[3800]  = 77;
  ram[3801]  = 77;
  ram[3802]  = 77;
  ram[3803]  = 77;
  ram[3804]  = 77;
  ram[3805]  = 76;
  ram[3806]  = 76;
  ram[3807]  = 76;
  ram[3808]  = 76;
  ram[3809]  = 76;
  ram[3810]  = 76;
  ram[3811]  = 75;
  ram[3812]  = 75;
  ram[3813]  = 75;
  ram[3814]  = 75;
  ram[3815]  = 75;
  ram[3816]  = 76;
  ram[3817]  = 76;
  ram[3818]  = 75;
  ram[3819]  = 75;
  ram[3820]  = 77;
  ram[3821]  = 77;
  ram[3822]  = 77;
  ram[3823]  = 77;
  ram[3824]  = 77;
  ram[3825]  = 77;
  ram[3826]  = 78;
  ram[3827]  = 76;
  ram[3828]  = 76;
  ram[3829]  = 76;
  ram[3830]  = 76;
  ram[3831]  = 76;
  ram[3832]  = 75;
  ram[3833]  = 75;
  ram[3834]  = 75;
  ram[3835]  = 75;
  ram[3836]  = 74;
  ram[3837]  = 73;
  ram[3838]  = 73;
  ram[3839]  = 72;
  ram[3840]  = 77;
  ram[3841]  = 77;
  ram[3842]  = 76;
  ram[3843]  = 75;
  ram[3844]  = 75;
  ram[3845]  = 75;
  ram[3846]  = 75;
  ram[3847]  = 75;
  ram[3848]  = 75;
  ram[3849]  = 75;
  ram[3850]  = 75;
  ram[3851]  = 75;
  ram[3852]  = 75;
  ram[3853]  = 75;
  ram[3854]  = 75;
  ram[3855]  = 75;
  ram[3856]  = 74;
  ram[3857]  = 74;
  ram[3858]  = 74;
  ram[3859]  = 74;
  ram[3860]  = 74;
  ram[3861]  = 74;
  ram[3862]  = 75;
  ram[3863]  = 75;
  ram[3864]  = 74;
  ram[3865]  = 74;
  ram[3866]  = 74;
  ram[3867]  = 74;
  ram[3868]  = 74;
  ram[3869]  = 74;
  ram[3870]  = 74;
  ram[3871]  = 74;
  ram[3872]  = 74;
  ram[3873]  = 74;
  ram[3874]  = 74;
  ram[3875]  = 74;
  ram[3876]  = 74;
  ram[3877]  = 74;
  ram[3878]  = 74;
  ram[3879]  = 74;
  ram[3880]  = 74;
  ram[3881]  = 74;
  ram[3882]  = 74;
  ram[3883]  = 74;
  ram[3884]  = 74;
  ram[3885]  = 74;
  ram[3886]  = 74;
  ram[3887]  = 74;
  ram[3888]  = 74;
  ram[3889]  = 74;
  ram[3890]  = 75;
  ram[3891]  = 74;
  ram[3892]  = 74;
  ram[3893]  = 74;
  ram[3894]  = 74;
  ram[3895]  = 75;
  ram[3896]  = 75;
  ram[3897]  = 75;
  ram[3898]  = 75;
  ram[3899]  = 75;
  ram[3900]  = 74;
  ram[3901]  = 74;
  ram[3902]  = 73;
  ram[3903]  = 72;
  ram[3904]  = 76;
  ram[3905]  = 77;
  ram[3906]  = 76;
  ram[3907]  = 75;
  ram[3908]  = 74;
  ram[3909]  = 75;
  ram[3910]  = 75;
  ram[3911]  = 74;
  ram[3912]  = 74;
  ram[3913]  = 74;
  ram[3914]  = 74;
  ram[3915]  = 74;
  ram[3916]  = 74;
  ram[3917]  = 74;
  ram[3918]  = 74;
  ram[3919]  = 74;
  ram[3920]  = 72;
  ram[3921]  = 72;
  ram[3922]  = 72;
  ram[3923]  = 73;
  ram[3924]  = 73;
  ram[3925]  = 73;
  ram[3926]  = 73;
  ram[3927]  = 73;
  ram[3928]  = 73;
  ram[3929]  = 72;
  ram[3930]  = 72;
  ram[3931]  = 72;
  ram[3932]  = 72;
  ram[3933]  = 72;
  ram[3934]  = 72;
  ram[3935]  = 72;
  ram[3936]  = 72;
  ram[3937]  = 72;
  ram[3938]  = 72;
  ram[3939]  = 72;
  ram[3940]  = 72;
  ram[3941]  = 72;
  ram[3942]  = 72;
  ram[3943]  = 72;
  ram[3944]  = 72;
  ram[3945]  = 72;
  ram[3946]  = 72;
  ram[3947]  = 72;
  ram[3948]  = 72;
  ram[3949]  = 72;
  ram[3950]  = 72;
  ram[3951]  = 72;
  ram[3952]  = 72;
  ram[3953]  = 72;
  ram[3954]  = 72;
  ram[3955]  = 72;
  ram[3956]  = 73;
  ram[3957]  = 73;
  ram[3958]  = 73;
  ram[3959]  = 73;
  ram[3960]  = 75;
  ram[3961]  = 75;
  ram[3962]  = 75;
  ram[3963]  = 75;
  ram[3964]  = 74;
  ram[3965]  = 74;
  ram[3966]  = 73;
  ram[3967]  = 72;
  ram[3968]  = 74;
  ram[3969]  = 75;
  ram[3970]  = 75;
  ram[3971]  = 74;
  ram[3972]  = 74;
  ram[3973]  = 75;
  ram[3974]  = 75;
  ram[3975]  = 75;
  ram[3976]  = 77;
  ram[3977]  = 77;
  ram[3978]  = 77;
  ram[3979]  = 77;
  ram[3980]  = 77;
  ram[3981]  = 77;
  ram[3982]  = 77;
  ram[3983]  = 77;
  ram[3984]  = 74;
  ram[3985]  = 74;
  ram[3986]  = 75;
  ram[3987]  = 75;
  ram[3988]  = 75;
  ram[3989]  = 75;
  ram[3990]  = 75;
  ram[3991]  = 75;
  ram[3992]  = 75;
  ram[3993]  = 75;
  ram[3994]  = 75;
  ram[3995]  = 75;
  ram[3996]  = 75;
  ram[3997]  = 75;
  ram[3998]  = 75;
  ram[3999]  = 75;
  ram[4000]  = 75;
  ram[4001]  = 75;
  ram[4002]  = 75;
  ram[4003]  = 75;
  ram[4004]  = 76;
  ram[4005]  = 76;
  ram[4006]  = 76;
  ram[4007]  = 76;
  ram[4008]  = 76;
  ram[4009]  = 76;
  ram[4010]  = 76;
  ram[4011]  = 76;
  ram[4012]  = 75;
  ram[4013]  = 75;
  ram[4014]  = 75;
  ram[4015]  = 75;
  ram[4016]  = 75;
  ram[4017]  = 75;
  ram[4018]  = 75;
  ram[4019]  = 75;
  ram[4020]  = 75;
  ram[4021]  = 75;
  ram[4022]  = 75;
  ram[4023]  = 75;
  ram[4024]  = 74;
  ram[4025]  = 74;
  ram[4026]  = 75;
  ram[4027]  = 75;
  ram[4028]  = 74;
  ram[4029]  = 74;
  ram[4030]  = 73;
  ram[4031]  = 72;
  ram[4032]  = 72;
  ram[4033]  = 73;
  ram[4034]  = 74;
  ram[4035]  = 74;
  ram[4036]  = 75;
  ram[4037]  = 76;
  ram[4038]  = 76;
  ram[4039]  = 75;
  ram[4040]  = 74;
  ram[4041]  = 74;
  ram[4042]  = 74;
  ram[4043]  = 74;
  ram[4044]  = 74;
  ram[4045]  = 74;
  ram[4046]  = 74;
  ram[4047]  = 74;
  ram[4048]  = 73;
  ram[4049]  = 73;
  ram[4050]  = 73;
  ram[4051]  = 73;
  ram[4052]  = 73;
  ram[4053]  = 73;
  ram[4054]  = 73;
  ram[4055]  = 73;
  ram[4056]  = 73;
  ram[4057]  = 73;
  ram[4058]  = 73;
  ram[4059]  = 73;
  ram[4060]  = 73;
  ram[4061]  = 73;
  ram[4062]  = 73;
  ram[4063]  = 73;
  ram[4064]  = 73;
  ram[4065]  = 73;
  ram[4066]  = 73;
  ram[4067]  = 73;
  ram[4068]  = 74;
  ram[4069]  = 74;
  ram[4070]  = 74;
  ram[4071]  = 74;
  ram[4072]  = 74;
  ram[4073]  = 74;
  ram[4074]  = 74;
  ram[4075]  = 74;
  ram[4076]  = 74;
  ram[4077]  = 74;
  ram[4078]  = 73;
  ram[4079]  = 73;
  ram[4080]  = 74;
  ram[4081]  = 74;
  ram[4082]  = 73;
  ram[4083]  = 73;
  ram[4084]  = 73;
  ram[4085]  = 74;
  ram[4086]  = 74;
  ram[4087]  = 74;
  ram[4088]  = 74;
  ram[4089]  = 74;
  ram[4090]  = 75;
  ram[4091]  = 75;
  ram[4092]  = 74;
  ram[4093]  = 74;
  ram[4094]  = 73;
  ram[4095]  = 72;
end

always @(posedge clock) begin
  dout <= ram[address];
end

endmodule
